-- megafunction wizard: %PARALLEL_ADD%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: parallel_add 

-- ============================================================
-- File Name: mapping_add.vhd
-- Megafunction Name(s):
-- 			parallel_add
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 15.0.0 Build 145 04/22/2015 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus II License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY mapping_add IS
	PORT
	(
		clock		: IN STD_LOGIC  := '0';
		data0x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data10x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data11x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data12x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data13x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data14x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data15x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data16x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data17x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data18x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data19x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data20x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data21x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data22x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data23x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data24x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data25x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data26x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data27x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data28x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data29x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data30x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data31x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data32x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data33x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data34x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data35x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data36x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data37x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data8x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		data9x		: IN STD_LOGIC_VECTOR (37 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (43 DOWNTO 0)
	);
END mapping_add;


ARCHITECTURE SYN OF mapping_add IS

--	type ALTERA_MF_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire1	: ALTERA_MF_LOGIC_2D (37 DOWNTO 0, 37 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire14	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire15	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire16	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire17	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire18	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire19	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire20	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire21	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire22	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire23	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire24	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire25	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire26	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire27	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire28	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire29	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire30	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire31	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire32	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire33	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire34	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire35	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire36	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire37	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire38	: STD_LOGIC_VECTOR (37 DOWNTO 0);
	SIGNAL sub_wire39	: STD_LOGIC_VECTOR (43 DOWNTO 0);

BEGIN
	sub_wire38    <= data0x(37 DOWNTO 0);
	sub_wire37    <= data1x(37 DOWNTO 0);
	sub_wire36    <= data2x(37 DOWNTO 0);
	sub_wire35    <= data3x(37 DOWNTO 0);
	sub_wire34    <= data4x(37 DOWNTO 0);
	sub_wire33    <= data5x(37 DOWNTO 0);
	sub_wire32    <= data6x(37 DOWNTO 0);
	sub_wire31    <= data7x(37 DOWNTO 0);
	sub_wire30    <= data8x(37 DOWNTO 0);
	sub_wire29    <= data9x(37 DOWNTO 0);
	sub_wire28    <= data10x(37 DOWNTO 0);
	sub_wire27    <= data11x(37 DOWNTO 0);
	sub_wire26    <= data12x(37 DOWNTO 0);
	sub_wire25    <= data13x(37 DOWNTO 0);
	sub_wire24    <= data14x(37 DOWNTO 0);
	sub_wire23    <= data15x(37 DOWNTO 0);
	sub_wire22    <= data16x(37 DOWNTO 0);
	sub_wire21    <= data17x(37 DOWNTO 0);
	sub_wire20    <= data18x(37 DOWNTO 0);
	sub_wire19    <= data19x(37 DOWNTO 0);
	sub_wire18    <= data20x(37 DOWNTO 0);
	sub_wire17    <= data21x(37 DOWNTO 0);
	sub_wire16    <= data22x(37 DOWNTO 0);
	sub_wire15    <= data23x(37 DOWNTO 0);
	sub_wire14    <= data24x(37 DOWNTO 0);
	sub_wire13    <= data25x(37 DOWNTO 0);
	sub_wire12    <= data26x(37 DOWNTO 0);
	sub_wire11    <= data27x(37 DOWNTO 0);
	sub_wire10    <= data28x(37 DOWNTO 0);
	sub_wire9    <= data29x(37 DOWNTO 0);
	sub_wire8    <= data30x(37 DOWNTO 0);
	sub_wire7    <= data31x(37 DOWNTO 0);
	sub_wire6    <= data32x(37 DOWNTO 0);
	sub_wire5    <= data33x(37 DOWNTO 0);
	sub_wire4    <= data34x(37 DOWNTO 0);
	sub_wire3    <= data35x(37 DOWNTO 0);
	sub_wire2    <= data36x(37 DOWNTO 0);
	sub_wire0    <= data37x(37 DOWNTO 0);
	sub_wire1(37, 0)    <= sub_wire0(0);
	sub_wire1(37, 1)    <= sub_wire0(1);
	sub_wire1(37, 2)    <= sub_wire0(2);
	sub_wire1(37, 3)    <= sub_wire0(3);
	sub_wire1(37, 4)    <= sub_wire0(4);
	sub_wire1(37, 5)    <= sub_wire0(5);
	sub_wire1(37, 6)    <= sub_wire0(6);
	sub_wire1(37, 7)    <= sub_wire0(7);
	sub_wire1(37, 8)    <= sub_wire0(8);
	sub_wire1(37, 9)    <= sub_wire0(9);
	sub_wire1(37, 10)    <= sub_wire0(10);
	sub_wire1(37, 11)    <= sub_wire0(11);
	sub_wire1(37, 12)    <= sub_wire0(12);
	sub_wire1(37, 13)    <= sub_wire0(13);
	sub_wire1(37, 14)    <= sub_wire0(14);
	sub_wire1(37, 15)    <= sub_wire0(15);
	sub_wire1(37, 16)    <= sub_wire0(16);
	sub_wire1(37, 17)    <= sub_wire0(17);
	sub_wire1(37, 18)    <= sub_wire0(18);
	sub_wire1(37, 19)    <= sub_wire0(19);
	sub_wire1(37, 20)    <= sub_wire0(20);
	sub_wire1(37, 21)    <= sub_wire0(21);
	sub_wire1(37, 22)    <= sub_wire0(22);
	sub_wire1(37, 23)    <= sub_wire0(23);
	sub_wire1(37, 24)    <= sub_wire0(24);
	sub_wire1(37, 25)    <= sub_wire0(25);
	sub_wire1(37, 26)    <= sub_wire0(26);
	sub_wire1(37, 27)    <= sub_wire0(27);
	sub_wire1(37, 28)    <= sub_wire0(28);
	sub_wire1(37, 29)    <= sub_wire0(29);
	sub_wire1(37, 30)    <= sub_wire0(30);
	sub_wire1(37, 31)    <= sub_wire0(31);
	sub_wire1(37, 32)    <= sub_wire0(32);
	sub_wire1(37, 33)    <= sub_wire0(33);
	sub_wire1(37, 34)    <= sub_wire0(34);
	sub_wire1(37, 35)    <= sub_wire0(35);
	sub_wire1(37, 36)    <= sub_wire0(36);
	sub_wire1(37, 37)    <= sub_wire0(37);
	sub_wire1(36, 0)    <= sub_wire2(0);
	sub_wire1(36, 1)    <= sub_wire2(1);
	sub_wire1(36, 2)    <= sub_wire2(2);
	sub_wire1(36, 3)    <= sub_wire2(3);
	sub_wire1(36, 4)    <= sub_wire2(4);
	sub_wire1(36, 5)    <= sub_wire2(5);
	sub_wire1(36, 6)    <= sub_wire2(6);
	sub_wire1(36, 7)    <= sub_wire2(7);
	sub_wire1(36, 8)    <= sub_wire2(8);
	sub_wire1(36, 9)    <= sub_wire2(9);
	sub_wire1(36, 10)    <= sub_wire2(10);
	sub_wire1(36, 11)    <= sub_wire2(11);
	sub_wire1(36, 12)    <= sub_wire2(12);
	sub_wire1(36, 13)    <= sub_wire2(13);
	sub_wire1(36, 14)    <= sub_wire2(14);
	sub_wire1(36, 15)    <= sub_wire2(15);
	sub_wire1(36, 16)    <= sub_wire2(16);
	sub_wire1(36, 17)    <= sub_wire2(17);
	sub_wire1(36, 18)    <= sub_wire2(18);
	sub_wire1(36, 19)    <= sub_wire2(19);
	sub_wire1(36, 20)    <= sub_wire2(20);
	sub_wire1(36, 21)    <= sub_wire2(21);
	sub_wire1(36, 22)    <= sub_wire2(22);
	sub_wire1(36, 23)    <= sub_wire2(23);
	sub_wire1(36, 24)    <= sub_wire2(24);
	sub_wire1(36, 25)    <= sub_wire2(25);
	sub_wire1(36, 26)    <= sub_wire2(26);
	sub_wire1(36, 27)    <= sub_wire2(27);
	sub_wire1(36, 28)    <= sub_wire2(28);
	sub_wire1(36, 29)    <= sub_wire2(29);
	sub_wire1(36, 30)    <= sub_wire2(30);
	sub_wire1(36, 31)    <= sub_wire2(31);
	sub_wire1(36, 32)    <= sub_wire2(32);
	sub_wire1(36, 33)    <= sub_wire2(33);
	sub_wire1(36, 34)    <= sub_wire2(34);
	sub_wire1(36, 35)    <= sub_wire2(35);
	sub_wire1(36, 36)    <= sub_wire2(36);
	sub_wire1(36, 37)    <= sub_wire2(37);
	sub_wire1(35, 0)    <= sub_wire3(0);
	sub_wire1(35, 1)    <= sub_wire3(1);
	sub_wire1(35, 2)    <= sub_wire3(2);
	sub_wire1(35, 3)    <= sub_wire3(3);
	sub_wire1(35, 4)    <= sub_wire3(4);
	sub_wire1(35, 5)    <= sub_wire3(5);
	sub_wire1(35, 6)    <= sub_wire3(6);
	sub_wire1(35, 7)    <= sub_wire3(7);
	sub_wire1(35, 8)    <= sub_wire3(8);
	sub_wire1(35, 9)    <= sub_wire3(9);
	sub_wire1(35, 10)    <= sub_wire3(10);
	sub_wire1(35, 11)    <= sub_wire3(11);
	sub_wire1(35, 12)    <= sub_wire3(12);
	sub_wire1(35, 13)    <= sub_wire3(13);
	sub_wire1(35, 14)    <= sub_wire3(14);
	sub_wire1(35, 15)    <= sub_wire3(15);
	sub_wire1(35, 16)    <= sub_wire3(16);
	sub_wire1(35, 17)    <= sub_wire3(17);
	sub_wire1(35, 18)    <= sub_wire3(18);
	sub_wire1(35, 19)    <= sub_wire3(19);
	sub_wire1(35, 20)    <= sub_wire3(20);
	sub_wire1(35, 21)    <= sub_wire3(21);
	sub_wire1(35, 22)    <= sub_wire3(22);
	sub_wire1(35, 23)    <= sub_wire3(23);
	sub_wire1(35, 24)    <= sub_wire3(24);
	sub_wire1(35, 25)    <= sub_wire3(25);
	sub_wire1(35, 26)    <= sub_wire3(26);
	sub_wire1(35, 27)    <= sub_wire3(27);
	sub_wire1(35, 28)    <= sub_wire3(28);
	sub_wire1(35, 29)    <= sub_wire3(29);
	sub_wire1(35, 30)    <= sub_wire3(30);
	sub_wire1(35, 31)    <= sub_wire3(31);
	sub_wire1(35, 32)    <= sub_wire3(32);
	sub_wire1(35, 33)    <= sub_wire3(33);
	sub_wire1(35, 34)    <= sub_wire3(34);
	sub_wire1(35, 35)    <= sub_wire3(35);
	sub_wire1(35, 36)    <= sub_wire3(36);
	sub_wire1(35, 37)    <= sub_wire3(37);
	sub_wire1(34, 0)    <= sub_wire4(0);
	sub_wire1(34, 1)    <= sub_wire4(1);
	sub_wire1(34, 2)    <= sub_wire4(2);
	sub_wire1(34, 3)    <= sub_wire4(3);
	sub_wire1(34, 4)    <= sub_wire4(4);
	sub_wire1(34, 5)    <= sub_wire4(5);
	sub_wire1(34, 6)    <= sub_wire4(6);
	sub_wire1(34, 7)    <= sub_wire4(7);
	sub_wire1(34, 8)    <= sub_wire4(8);
	sub_wire1(34, 9)    <= sub_wire4(9);
	sub_wire1(34, 10)    <= sub_wire4(10);
	sub_wire1(34, 11)    <= sub_wire4(11);
	sub_wire1(34, 12)    <= sub_wire4(12);
	sub_wire1(34, 13)    <= sub_wire4(13);
	sub_wire1(34, 14)    <= sub_wire4(14);
	sub_wire1(34, 15)    <= sub_wire4(15);
	sub_wire1(34, 16)    <= sub_wire4(16);
	sub_wire1(34, 17)    <= sub_wire4(17);
	sub_wire1(34, 18)    <= sub_wire4(18);
	sub_wire1(34, 19)    <= sub_wire4(19);
	sub_wire1(34, 20)    <= sub_wire4(20);
	sub_wire1(34, 21)    <= sub_wire4(21);
	sub_wire1(34, 22)    <= sub_wire4(22);
	sub_wire1(34, 23)    <= sub_wire4(23);
	sub_wire1(34, 24)    <= sub_wire4(24);
	sub_wire1(34, 25)    <= sub_wire4(25);
	sub_wire1(34, 26)    <= sub_wire4(26);
	sub_wire1(34, 27)    <= sub_wire4(27);
	sub_wire1(34, 28)    <= sub_wire4(28);
	sub_wire1(34, 29)    <= sub_wire4(29);
	sub_wire1(34, 30)    <= sub_wire4(30);
	sub_wire1(34, 31)    <= sub_wire4(31);
	sub_wire1(34, 32)    <= sub_wire4(32);
	sub_wire1(34, 33)    <= sub_wire4(33);
	sub_wire1(34, 34)    <= sub_wire4(34);
	sub_wire1(34, 35)    <= sub_wire4(35);
	sub_wire1(34, 36)    <= sub_wire4(36);
	sub_wire1(34, 37)    <= sub_wire4(37);
	sub_wire1(33, 0)    <= sub_wire5(0);
	sub_wire1(33, 1)    <= sub_wire5(1);
	sub_wire1(33, 2)    <= sub_wire5(2);
	sub_wire1(33, 3)    <= sub_wire5(3);
	sub_wire1(33, 4)    <= sub_wire5(4);
	sub_wire1(33, 5)    <= sub_wire5(5);
	sub_wire1(33, 6)    <= sub_wire5(6);
	sub_wire1(33, 7)    <= sub_wire5(7);
	sub_wire1(33, 8)    <= sub_wire5(8);
	sub_wire1(33, 9)    <= sub_wire5(9);
	sub_wire1(33, 10)    <= sub_wire5(10);
	sub_wire1(33, 11)    <= sub_wire5(11);
	sub_wire1(33, 12)    <= sub_wire5(12);
	sub_wire1(33, 13)    <= sub_wire5(13);
	sub_wire1(33, 14)    <= sub_wire5(14);
	sub_wire1(33, 15)    <= sub_wire5(15);
	sub_wire1(33, 16)    <= sub_wire5(16);
	sub_wire1(33, 17)    <= sub_wire5(17);
	sub_wire1(33, 18)    <= sub_wire5(18);
	sub_wire1(33, 19)    <= sub_wire5(19);
	sub_wire1(33, 20)    <= sub_wire5(20);
	sub_wire1(33, 21)    <= sub_wire5(21);
	sub_wire1(33, 22)    <= sub_wire5(22);
	sub_wire1(33, 23)    <= sub_wire5(23);
	sub_wire1(33, 24)    <= sub_wire5(24);
	sub_wire1(33, 25)    <= sub_wire5(25);
	sub_wire1(33, 26)    <= sub_wire5(26);
	sub_wire1(33, 27)    <= sub_wire5(27);
	sub_wire1(33, 28)    <= sub_wire5(28);
	sub_wire1(33, 29)    <= sub_wire5(29);
	sub_wire1(33, 30)    <= sub_wire5(30);
	sub_wire1(33, 31)    <= sub_wire5(31);
	sub_wire1(33, 32)    <= sub_wire5(32);
	sub_wire1(33, 33)    <= sub_wire5(33);
	sub_wire1(33, 34)    <= sub_wire5(34);
	sub_wire1(33, 35)    <= sub_wire5(35);
	sub_wire1(33, 36)    <= sub_wire5(36);
	sub_wire1(33, 37)    <= sub_wire5(37);
	sub_wire1(32, 0)    <= sub_wire6(0);
	sub_wire1(32, 1)    <= sub_wire6(1);
	sub_wire1(32, 2)    <= sub_wire6(2);
	sub_wire1(32, 3)    <= sub_wire6(3);
	sub_wire1(32, 4)    <= sub_wire6(4);
	sub_wire1(32, 5)    <= sub_wire6(5);
	sub_wire1(32, 6)    <= sub_wire6(6);
	sub_wire1(32, 7)    <= sub_wire6(7);
	sub_wire1(32, 8)    <= sub_wire6(8);
	sub_wire1(32, 9)    <= sub_wire6(9);
	sub_wire1(32, 10)    <= sub_wire6(10);
	sub_wire1(32, 11)    <= sub_wire6(11);
	sub_wire1(32, 12)    <= sub_wire6(12);
	sub_wire1(32, 13)    <= sub_wire6(13);
	sub_wire1(32, 14)    <= sub_wire6(14);
	sub_wire1(32, 15)    <= sub_wire6(15);
	sub_wire1(32, 16)    <= sub_wire6(16);
	sub_wire1(32, 17)    <= sub_wire6(17);
	sub_wire1(32, 18)    <= sub_wire6(18);
	sub_wire1(32, 19)    <= sub_wire6(19);
	sub_wire1(32, 20)    <= sub_wire6(20);
	sub_wire1(32, 21)    <= sub_wire6(21);
	sub_wire1(32, 22)    <= sub_wire6(22);
	sub_wire1(32, 23)    <= sub_wire6(23);
	sub_wire1(32, 24)    <= sub_wire6(24);
	sub_wire1(32, 25)    <= sub_wire6(25);
	sub_wire1(32, 26)    <= sub_wire6(26);
	sub_wire1(32, 27)    <= sub_wire6(27);
	sub_wire1(32, 28)    <= sub_wire6(28);
	sub_wire1(32, 29)    <= sub_wire6(29);
	sub_wire1(32, 30)    <= sub_wire6(30);
	sub_wire1(32, 31)    <= sub_wire6(31);
	sub_wire1(32, 32)    <= sub_wire6(32);
	sub_wire1(32, 33)    <= sub_wire6(33);
	sub_wire1(32, 34)    <= sub_wire6(34);
	sub_wire1(32, 35)    <= sub_wire6(35);
	sub_wire1(32, 36)    <= sub_wire6(36);
	sub_wire1(32, 37)    <= sub_wire6(37);
	sub_wire1(31, 0)    <= sub_wire7(0);
	sub_wire1(31, 1)    <= sub_wire7(1);
	sub_wire1(31, 2)    <= sub_wire7(2);
	sub_wire1(31, 3)    <= sub_wire7(3);
	sub_wire1(31, 4)    <= sub_wire7(4);
	sub_wire1(31, 5)    <= sub_wire7(5);
	sub_wire1(31, 6)    <= sub_wire7(6);
	sub_wire1(31, 7)    <= sub_wire7(7);
	sub_wire1(31, 8)    <= sub_wire7(8);
	sub_wire1(31, 9)    <= sub_wire7(9);
	sub_wire1(31, 10)    <= sub_wire7(10);
	sub_wire1(31, 11)    <= sub_wire7(11);
	sub_wire1(31, 12)    <= sub_wire7(12);
	sub_wire1(31, 13)    <= sub_wire7(13);
	sub_wire1(31, 14)    <= sub_wire7(14);
	sub_wire1(31, 15)    <= sub_wire7(15);
	sub_wire1(31, 16)    <= sub_wire7(16);
	sub_wire1(31, 17)    <= sub_wire7(17);
	sub_wire1(31, 18)    <= sub_wire7(18);
	sub_wire1(31, 19)    <= sub_wire7(19);
	sub_wire1(31, 20)    <= sub_wire7(20);
	sub_wire1(31, 21)    <= sub_wire7(21);
	sub_wire1(31, 22)    <= sub_wire7(22);
	sub_wire1(31, 23)    <= sub_wire7(23);
	sub_wire1(31, 24)    <= sub_wire7(24);
	sub_wire1(31, 25)    <= sub_wire7(25);
	sub_wire1(31, 26)    <= sub_wire7(26);
	sub_wire1(31, 27)    <= sub_wire7(27);
	sub_wire1(31, 28)    <= sub_wire7(28);
	sub_wire1(31, 29)    <= sub_wire7(29);
	sub_wire1(31, 30)    <= sub_wire7(30);
	sub_wire1(31, 31)    <= sub_wire7(31);
	sub_wire1(31, 32)    <= sub_wire7(32);
	sub_wire1(31, 33)    <= sub_wire7(33);
	sub_wire1(31, 34)    <= sub_wire7(34);
	sub_wire1(31, 35)    <= sub_wire7(35);
	sub_wire1(31, 36)    <= sub_wire7(36);
	sub_wire1(31, 37)    <= sub_wire7(37);
	sub_wire1(30, 0)    <= sub_wire8(0);
	sub_wire1(30, 1)    <= sub_wire8(1);
	sub_wire1(30, 2)    <= sub_wire8(2);
	sub_wire1(30, 3)    <= sub_wire8(3);
	sub_wire1(30, 4)    <= sub_wire8(4);
	sub_wire1(30, 5)    <= sub_wire8(5);
	sub_wire1(30, 6)    <= sub_wire8(6);
	sub_wire1(30, 7)    <= sub_wire8(7);
	sub_wire1(30, 8)    <= sub_wire8(8);
	sub_wire1(30, 9)    <= sub_wire8(9);
	sub_wire1(30, 10)    <= sub_wire8(10);
	sub_wire1(30, 11)    <= sub_wire8(11);
	sub_wire1(30, 12)    <= sub_wire8(12);
	sub_wire1(30, 13)    <= sub_wire8(13);
	sub_wire1(30, 14)    <= sub_wire8(14);
	sub_wire1(30, 15)    <= sub_wire8(15);
	sub_wire1(30, 16)    <= sub_wire8(16);
	sub_wire1(30, 17)    <= sub_wire8(17);
	sub_wire1(30, 18)    <= sub_wire8(18);
	sub_wire1(30, 19)    <= sub_wire8(19);
	sub_wire1(30, 20)    <= sub_wire8(20);
	sub_wire1(30, 21)    <= sub_wire8(21);
	sub_wire1(30, 22)    <= sub_wire8(22);
	sub_wire1(30, 23)    <= sub_wire8(23);
	sub_wire1(30, 24)    <= sub_wire8(24);
	sub_wire1(30, 25)    <= sub_wire8(25);
	sub_wire1(30, 26)    <= sub_wire8(26);
	sub_wire1(30, 27)    <= sub_wire8(27);
	sub_wire1(30, 28)    <= sub_wire8(28);
	sub_wire1(30, 29)    <= sub_wire8(29);
	sub_wire1(30, 30)    <= sub_wire8(30);
	sub_wire1(30, 31)    <= sub_wire8(31);
	sub_wire1(30, 32)    <= sub_wire8(32);
	sub_wire1(30, 33)    <= sub_wire8(33);
	sub_wire1(30, 34)    <= sub_wire8(34);
	sub_wire1(30, 35)    <= sub_wire8(35);
	sub_wire1(30, 36)    <= sub_wire8(36);
	sub_wire1(30, 37)    <= sub_wire8(37);
	sub_wire1(29, 0)    <= sub_wire9(0);
	sub_wire1(29, 1)    <= sub_wire9(1);
	sub_wire1(29, 2)    <= sub_wire9(2);
	sub_wire1(29, 3)    <= sub_wire9(3);
	sub_wire1(29, 4)    <= sub_wire9(4);
	sub_wire1(29, 5)    <= sub_wire9(5);
	sub_wire1(29, 6)    <= sub_wire9(6);
	sub_wire1(29, 7)    <= sub_wire9(7);
	sub_wire1(29, 8)    <= sub_wire9(8);
	sub_wire1(29, 9)    <= sub_wire9(9);
	sub_wire1(29, 10)    <= sub_wire9(10);
	sub_wire1(29, 11)    <= sub_wire9(11);
	sub_wire1(29, 12)    <= sub_wire9(12);
	sub_wire1(29, 13)    <= sub_wire9(13);
	sub_wire1(29, 14)    <= sub_wire9(14);
	sub_wire1(29, 15)    <= sub_wire9(15);
	sub_wire1(29, 16)    <= sub_wire9(16);
	sub_wire1(29, 17)    <= sub_wire9(17);
	sub_wire1(29, 18)    <= sub_wire9(18);
	sub_wire1(29, 19)    <= sub_wire9(19);
	sub_wire1(29, 20)    <= sub_wire9(20);
	sub_wire1(29, 21)    <= sub_wire9(21);
	sub_wire1(29, 22)    <= sub_wire9(22);
	sub_wire1(29, 23)    <= sub_wire9(23);
	sub_wire1(29, 24)    <= sub_wire9(24);
	sub_wire1(29, 25)    <= sub_wire9(25);
	sub_wire1(29, 26)    <= sub_wire9(26);
	sub_wire1(29, 27)    <= sub_wire9(27);
	sub_wire1(29, 28)    <= sub_wire9(28);
	sub_wire1(29, 29)    <= sub_wire9(29);
	sub_wire1(29, 30)    <= sub_wire9(30);
	sub_wire1(29, 31)    <= sub_wire9(31);
	sub_wire1(29, 32)    <= sub_wire9(32);
	sub_wire1(29, 33)    <= sub_wire9(33);
	sub_wire1(29, 34)    <= sub_wire9(34);
	sub_wire1(29, 35)    <= sub_wire9(35);
	sub_wire1(29, 36)    <= sub_wire9(36);
	sub_wire1(29, 37)    <= sub_wire9(37);
	sub_wire1(28, 0)    <= sub_wire10(0);
	sub_wire1(28, 1)    <= sub_wire10(1);
	sub_wire1(28, 2)    <= sub_wire10(2);
	sub_wire1(28, 3)    <= sub_wire10(3);
	sub_wire1(28, 4)    <= sub_wire10(4);
	sub_wire1(28, 5)    <= sub_wire10(5);
	sub_wire1(28, 6)    <= sub_wire10(6);
	sub_wire1(28, 7)    <= sub_wire10(7);
	sub_wire1(28, 8)    <= sub_wire10(8);
	sub_wire1(28, 9)    <= sub_wire10(9);
	sub_wire1(28, 10)    <= sub_wire10(10);
	sub_wire1(28, 11)    <= sub_wire10(11);
	sub_wire1(28, 12)    <= sub_wire10(12);
	sub_wire1(28, 13)    <= sub_wire10(13);
	sub_wire1(28, 14)    <= sub_wire10(14);
	sub_wire1(28, 15)    <= sub_wire10(15);
	sub_wire1(28, 16)    <= sub_wire10(16);
	sub_wire1(28, 17)    <= sub_wire10(17);
	sub_wire1(28, 18)    <= sub_wire10(18);
	sub_wire1(28, 19)    <= sub_wire10(19);
	sub_wire1(28, 20)    <= sub_wire10(20);
	sub_wire1(28, 21)    <= sub_wire10(21);
	sub_wire1(28, 22)    <= sub_wire10(22);
	sub_wire1(28, 23)    <= sub_wire10(23);
	sub_wire1(28, 24)    <= sub_wire10(24);
	sub_wire1(28, 25)    <= sub_wire10(25);
	sub_wire1(28, 26)    <= sub_wire10(26);
	sub_wire1(28, 27)    <= sub_wire10(27);
	sub_wire1(28, 28)    <= sub_wire10(28);
	sub_wire1(28, 29)    <= sub_wire10(29);
	sub_wire1(28, 30)    <= sub_wire10(30);
	sub_wire1(28, 31)    <= sub_wire10(31);
	sub_wire1(28, 32)    <= sub_wire10(32);
	sub_wire1(28, 33)    <= sub_wire10(33);
	sub_wire1(28, 34)    <= sub_wire10(34);
	sub_wire1(28, 35)    <= sub_wire10(35);
	sub_wire1(28, 36)    <= sub_wire10(36);
	sub_wire1(28, 37)    <= sub_wire10(37);
	sub_wire1(27, 0)    <= sub_wire11(0);
	sub_wire1(27, 1)    <= sub_wire11(1);
	sub_wire1(27, 2)    <= sub_wire11(2);
	sub_wire1(27, 3)    <= sub_wire11(3);
	sub_wire1(27, 4)    <= sub_wire11(4);
	sub_wire1(27, 5)    <= sub_wire11(5);
	sub_wire1(27, 6)    <= sub_wire11(6);
	sub_wire1(27, 7)    <= sub_wire11(7);
	sub_wire1(27, 8)    <= sub_wire11(8);
	sub_wire1(27, 9)    <= sub_wire11(9);
	sub_wire1(27, 10)    <= sub_wire11(10);
	sub_wire1(27, 11)    <= sub_wire11(11);
	sub_wire1(27, 12)    <= sub_wire11(12);
	sub_wire1(27, 13)    <= sub_wire11(13);
	sub_wire1(27, 14)    <= sub_wire11(14);
	sub_wire1(27, 15)    <= sub_wire11(15);
	sub_wire1(27, 16)    <= sub_wire11(16);
	sub_wire1(27, 17)    <= sub_wire11(17);
	sub_wire1(27, 18)    <= sub_wire11(18);
	sub_wire1(27, 19)    <= sub_wire11(19);
	sub_wire1(27, 20)    <= sub_wire11(20);
	sub_wire1(27, 21)    <= sub_wire11(21);
	sub_wire1(27, 22)    <= sub_wire11(22);
	sub_wire1(27, 23)    <= sub_wire11(23);
	sub_wire1(27, 24)    <= sub_wire11(24);
	sub_wire1(27, 25)    <= sub_wire11(25);
	sub_wire1(27, 26)    <= sub_wire11(26);
	sub_wire1(27, 27)    <= sub_wire11(27);
	sub_wire1(27, 28)    <= sub_wire11(28);
	sub_wire1(27, 29)    <= sub_wire11(29);
	sub_wire1(27, 30)    <= sub_wire11(30);
	sub_wire1(27, 31)    <= sub_wire11(31);
	sub_wire1(27, 32)    <= sub_wire11(32);
	sub_wire1(27, 33)    <= sub_wire11(33);
	sub_wire1(27, 34)    <= sub_wire11(34);
	sub_wire1(27, 35)    <= sub_wire11(35);
	sub_wire1(27, 36)    <= sub_wire11(36);
	sub_wire1(27, 37)    <= sub_wire11(37);
	sub_wire1(26, 0)    <= sub_wire12(0);
	sub_wire1(26, 1)    <= sub_wire12(1);
	sub_wire1(26, 2)    <= sub_wire12(2);
	sub_wire1(26, 3)    <= sub_wire12(3);
	sub_wire1(26, 4)    <= sub_wire12(4);
	sub_wire1(26, 5)    <= sub_wire12(5);
	sub_wire1(26, 6)    <= sub_wire12(6);
	sub_wire1(26, 7)    <= sub_wire12(7);
	sub_wire1(26, 8)    <= sub_wire12(8);
	sub_wire1(26, 9)    <= sub_wire12(9);
	sub_wire1(26, 10)    <= sub_wire12(10);
	sub_wire1(26, 11)    <= sub_wire12(11);
	sub_wire1(26, 12)    <= sub_wire12(12);
	sub_wire1(26, 13)    <= sub_wire12(13);
	sub_wire1(26, 14)    <= sub_wire12(14);
	sub_wire1(26, 15)    <= sub_wire12(15);
	sub_wire1(26, 16)    <= sub_wire12(16);
	sub_wire1(26, 17)    <= sub_wire12(17);
	sub_wire1(26, 18)    <= sub_wire12(18);
	sub_wire1(26, 19)    <= sub_wire12(19);
	sub_wire1(26, 20)    <= sub_wire12(20);
	sub_wire1(26, 21)    <= sub_wire12(21);
	sub_wire1(26, 22)    <= sub_wire12(22);
	sub_wire1(26, 23)    <= sub_wire12(23);
	sub_wire1(26, 24)    <= sub_wire12(24);
	sub_wire1(26, 25)    <= sub_wire12(25);
	sub_wire1(26, 26)    <= sub_wire12(26);
	sub_wire1(26, 27)    <= sub_wire12(27);
	sub_wire1(26, 28)    <= sub_wire12(28);
	sub_wire1(26, 29)    <= sub_wire12(29);
	sub_wire1(26, 30)    <= sub_wire12(30);
	sub_wire1(26, 31)    <= sub_wire12(31);
	sub_wire1(26, 32)    <= sub_wire12(32);
	sub_wire1(26, 33)    <= sub_wire12(33);
	sub_wire1(26, 34)    <= sub_wire12(34);
	sub_wire1(26, 35)    <= sub_wire12(35);
	sub_wire1(26, 36)    <= sub_wire12(36);
	sub_wire1(26, 37)    <= sub_wire12(37);
	sub_wire1(25, 0)    <= sub_wire13(0);
	sub_wire1(25, 1)    <= sub_wire13(1);
	sub_wire1(25, 2)    <= sub_wire13(2);
	sub_wire1(25, 3)    <= sub_wire13(3);
	sub_wire1(25, 4)    <= sub_wire13(4);
	sub_wire1(25, 5)    <= sub_wire13(5);
	sub_wire1(25, 6)    <= sub_wire13(6);
	sub_wire1(25, 7)    <= sub_wire13(7);
	sub_wire1(25, 8)    <= sub_wire13(8);
	sub_wire1(25, 9)    <= sub_wire13(9);
	sub_wire1(25, 10)    <= sub_wire13(10);
	sub_wire1(25, 11)    <= sub_wire13(11);
	sub_wire1(25, 12)    <= sub_wire13(12);
	sub_wire1(25, 13)    <= sub_wire13(13);
	sub_wire1(25, 14)    <= sub_wire13(14);
	sub_wire1(25, 15)    <= sub_wire13(15);
	sub_wire1(25, 16)    <= sub_wire13(16);
	sub_wire1(25, 17)    <= sub_wire13(17);
	sub_wire1(25, 18)    <= sub_wire13(18);
	sub_wire1(25, 19)    <= sub_wire13(19);
	sub_wire1(25, 20)    <= sub_wire13(20);
	sub_wire1(25, 21)    <= sub_wire13(21);
	sub_wire1(25, 22)    <= sub_wire13(22);
	sub_wire1(25, 23)    <= sub_wire13(23);
	sub_wire1(25, 24)    <= sub_wire13(24);
	sub_wire1(25, 25)    <= sub_wire13(25);
	sub_wire1(25, 26)    <= sub_wire13(26);
	sub_wire1(25, 27)    <= sub_wire13(27);
	sub_wire1(25, 28)    <= sub_wire13(28);
	sub_wire1(25, 29)    <= sub_wire13(29);
	sub_wire1(25, 30)    <= sub_wire13(30);
	sub_wire1(25, 31)    <= sub_wire13(31);
	sub_wire1(25, 32)    <= sub_wire13(32);
	sub_wire1(25, 33)    <= sub_wire13(33);
	sub_wire1(25, 34)    <= sub_wire13(34);
	sub_wire1(25, 35)    <= sub_wire13(35);
	sub_wire1(25, 36)    <= sub_wire13(36);
	sub_wire1(25, 37)    <= sub_wire13(37);
	sub_wire1(24, 0)    <= sub_wire14(0);
	sub_wire1(24, 1)    <= sub_wire14(1);
	sub_wire1(24, 2)    <= sub_wire14(2);
	sub_wire1(24, 3)    <= sub_wire14(3);
	sub_wire1(24, 4)    <= sub_wire14(4);
	sub_wire1(24, 5)    <= sub_wire14(5);
	sub_wire1(24, 6)    <= sub_wire14(6);
	sub_wire1(24, 7)    <= sub_wire14(7);
	sub_wire1(24, 8)    <= sub_wire14(8);
	sub_wire1(24, 9)    <= sub_wire14(9);
	sub_wire1(24, 10)    <= sub_wire14(10);
	sub_wire1(24, 11)    <= sub_wire14(11);
	sub_wire1(24, 12)    <= sub_wire14(12);
	sub_wire1(24, 13)    <= sub_wire14(13);
	sub_wire1(24, 14)    <= sub_wire14(14);
	sub_wire1(24, 15)    <= sub_wire14(15);
	sub_wire1(24, 16)    <= sub_wire14(16);
	sub_wire1(24, 17)    <= sub_wire14(17);
	sub_wire1(24, 18)    <= sub_wire14(18);
	sub_wire1(24, 19)    <= sub_wire14(19);
	sub_wire1(24, 20)    <= sub_wire14(20);
	sub_wire1(24, 21)    <= sub_wire14(21);
	sub_wire1(24, 22)    <= sub_wire14(22);
	sub_wire1(24, 23)    <= sub_wire14(23);
	sub_wire1(24, 24)    <= sub_wire14(24);
	sub_wire1(24, 25)    <= sub_wire14(25);
	sub_wire1(24, 26)    <= sub_wire14(26);
	sub_wire1(24, 27)    <= sub_wire14(27);
	sub_wire1(24, 28)    <= sub_wire14(28);
	sub_wire1(24, 29)    <= sub_wire14(29);
	sub_wire1(24, 30)    <= sub_wire14(30);
	sub_wire1(24, 31)    <= sub_wire14(31);
	sub_wire1(24, 32)    <= sub_wire14(32);
	sub_wire1(24, 33)    <= sub_wire14(33);
	sub_wire1(24, 34)    <= sub_wire14(34);
	sub_wire1(24, 35)    <= sub_wire14(35);
	sub_wire1(24, 36)    <= sub_wire14(36);
	sub_wire1(24, 37)    <= sub_wire14(37);
	sub_wire1(23, 0)    <= sub_wire15(0);
	sub_wire1(23, 1)    <= sub_wire15(1);
	sub_wire1(23, 2)    <= sub_wire15(2);
	sub_wire1(23, 3)    <= sub_wire15(3);
	sub_wire1(23, 4)    <= sub_wire15(4);
	sub_wire1(23, 5)    <= sub_wire15(5);
	sub_wire1(23, 6)    <= sub_wire15(6);
	sub_wire1(23, 7)    <= sub_wire15(7);
	sub_wire1(23, 8)    <= sub_wire15(8);
	sub_wire1(23, 9)    <= sub_wire15(9);
	sub_wire1(23, 10)    <= sub_wire15(10);
	sub_wire1(23, 11)    <= sub_wire15(11);
	sub_wire1(23, 12)    <= sub_wire15(12);
	sub_wire1(23, 13)    <= sub_wire15(13);
	sub_wire1(23, 14)    <= sub_wire15(14);
	sub_wire1(23, 15)    <= sub_wire15(15);
	sub_wire1(23, 16)    <= sub_wire15(16);
	sub_wire1(23, 17)    <= sub_wire15(17);
	sub_wire1(23, 18)    <= sub_wire15(18);
	sub_wire1(23, 19)    <= sub_wire15(19);
	sub_wire1(23, 20)    <= sub_wire15(20);
	sub_wire1(23, 21)    <= sub_wire15(21);
	sub_wire1(23, 22)    <= sub_wire15(22);
	sub_wire1(23, 23)    <= sub_wire15(23);
	sub_wire1(23, 24)    <= sub_wire15(24);
	sub_wire1(23, 25)    <= sub_wire15(25);
	sub_wire1(23, 26)    <= sub_wire15(26);
	sub_wire1(23, 27)    <= sub_wire15(27);
	sub_wire1(23, 28)    <= sub_wire15(28);
	sub_wire1(23, 29)    <= sub_wire15(29);
	sub_wire1(23, 30)    <= sub_wire15(30);
	sub_wire1(23, 31)    <= sub_wire15(31);
	sub_wire1(23, 32)    <= sub_wire15(32);
	sub_wire1(23, 33)    <= sub_wire15(33);
	sub_wire1(23, 34)    <= sub_wire15(34);
	sub_wire1(23, 35)    <= sub_wire15(35);
	sub_wire1(23, 36)    <= sub_wire15(36);
	sub_wire1(23, 37)    <= sub_wire15(37);
	sub_wire1(22, 0)    <= sub_wire16(0);
	sub_wire1(22, 1)    <= sub_wire16(1);
	sub_wire1(22, 2)    <= sub_wire16(2);
	sub_wire1(22, 3)    <= sub_wire16(3);
	sub_wire1(22, 4)    <= sub_wire16(4);
	sub_wire1(22, 5)    <= sub_wire16(5);
	sub_wire1(22, 6)    <= sub_wire16(6);
	sub_wire1(22, 7)    <= sub_wire16(7);
	sub_wire1(22, 8)    <= sub_wire16(8);
	sub_wire1(22, 9)    <= sub_wire16(9);
	sub_wire1(22, 10)    <= sub_wire16(10);
	sub_wire1(22, 11)    <= sub_wire16(11);
	sub_wire1(22, 12)    <= sub_wire16(12);
	sub_wire1(22, 13)    <= sub_wire16(13);
	sub_wire1(22, 14)    <= sub_wire16(14);
	sub_wire1(22, 15)    <= sub_wire16(15);
	sub_wire1(22, 16)    <= sub_wire16(16);
	sub_wire1(22, 17)    <= sub_wire16(17);
	sub_wire1(22, 18)    <= sub_wire16(18);
	sub_wire1(22, 19)    <= sub_wire16(19);
	sub_wire1(22, 20)    <= sub_wire16(20);
	sub_wire1(22, 21)    <= sub_wire16(21);
	sub_wire1(22, 22)    <= sub_wire16(22);
	sub_wire1(22, 23)    <= sub_wire16(23);
	sub_wire1(22, 24)    <= sub_wire16(24);
	sub_wire1(22, 25)    <= sub_wire16(25);
	sub_wire1(22, 26)    <= sub_wire16(26);
	sub_wire1(22, 27)    <= sub_wire16(27);
	sub_wire1(22, 28)    <= sub_wire16(28);
	sub_wire1(22, 29)    <= sub_wire16(29);
	sub_wire1(22, 30)    <= sub_wire16(30);
	sub_wire1(22, 31)    <= sub_wire16(31);
	sub_wire1(22, 32)    <= sub_wire16(32);
	sub_wire1(22, 33)    <= sub_wire16(33);
	sub_wire1(22, 34)    <= sub_wire16(34);
	sub_wire1(22, 35)    <= sub_wire16(35);
	sub_wire1(22, 36)    <= sub_wire16(36);
	sub_wire1(22, 37)    <= sub_wire16(37);
	sub_wire1(21, 0)    <= sub_wire17(0);
	sub_wire1(21, 1)    <= sub_wire17(1);
	sub_wire1(21, 2)    <= sub_wire17(2);
	sub_wire1(21, 3)    <= sub_wire17(3);
	sub_wire1(21, 4)    <= sub_wire17(4);
	sub_wire1(21, 5)    <= sub_wire17(5);
	sub_wire1(21, 6)    <= sub_wire17(6);
	sub_wire1(21, 7)    <= sub_wire17(7);
	sub_wire1(21, 8)    <= sub_wire17(8);
	sub_wire1(21, 9)    <= sub_wire17(9);
	sub_wire1(21, 10)    <= sub_wire17(10);
	sub_wire1(21, 11)    <= sub_wire17(11);
	sub_wire1(21, 12)    <= sub_wire17(12);
	sub_wire1(21, 13)    <= sub_wire17(13);
	sub_wire1(21, 14)    <= sub_wire17(14);
	sub_wire1(21, 15)    <= sub_wire17(15);
	sub_wire1(21, 16)    <= sub_wire17(16);
	sub_wire1(21, 17)    <= sub_wire17(17);
	sub_wire1(21, 18)    <= sub_wire17(18);
	sub_wire1(21, 19)    <= sub_wire17(19);
	sub_wire1(21, 20)    <= sub_wire17(20);
	sub_wire1(21, 21)    <= sub_wire17(21);
	sub_wire1(21, 22)    <= sub_wire17(22);
	sub_wire1(21, 23)    <= sub_wire17(23);
	sub_wire1(21, 24)    <= sub_wire17(24);
	sub_wire1(21, 25)    <= sub_wire17(25);
	sub_wire1(21, 26)    <= sub_wire17(26);
	sub_wire1(21, 27)    <= sub_wire17(27);
	sub_wire1(21, 28)    <= sub_wire17(28);
	sub_wire1(21, 29)    <= sub_wire17(29);
	sub_wire1(21, 30)    <= sub_wire17(30);
	sub_wire1(21, 31)    <= sub_wire17(31);
	sub_wire1(21, 32)    <= sub_wire17(32);
	sub_wire1(21, 33)    <= sub_wire17(33);
	sub_wire1(21, 34)    <= sub_wire17(34);
	sub_wire1(21, 35)    <= sub_wire17(35);
	sub_wire1(21, 36)    <= sub_wire17(36);
	sub_wire1(21, 37)    <= sub_wire17(37);
	sub_wire1(20, 0)    <= sub_wire18(0);
	sub_wire1(20, 1)    <= sub_wire18(1);
	sub_wire1(20, 2)    <= sub_wire18(2);
	sub_wire1(20, 3)    <= sub_wire18(3);
	sub_wire1(20, 4)    <= sub_wire18(4);
	sub_wire1(20, 5)    <= sub_wire18(5);
	sub_wire1(20, 6)    <= sub_wire18(6);
	sub_wire1(20, 7)    <= sub_wire18(7);
	sub_wire1(20, 8)    <= sub_wire18(8);
	sub_wire1(20, 9)    <= sub_wire18(9);
	sub_wire1(20, 10)    <= sub_wire18(10);
	sub_wire1(20, 11)    <= sub_wire18(11);
	sub_wire1(20, 12)    <= sub_wire18(12);
	sub_wire1(20, 13)    <= sub_wire18(13);
	sub_wire1(20, 14)    <= sub_wire18(14);
	sub_wire1(20, 15)    <= sub_wire18(15);
	sub_wire1(20, 16)    <= sub_wire18(16);
	sub_wire1(20, 17)    <= sub_wire18(17);
	sub_wire1(20, 18)    <= sub_wire18(18);
	sub_wire1(20, 19)    <= sub_wire18(19);
	sub_wire1(20, 20)    <= sub_wire18(20);
	sub_wire1(20, 21)    <= sub_wire18(21);
	sub_wire1(20, 22)    <= sub_wire18(22);
	sub_wire1(20, 23)    <= sub_wire18(23);
	sub_wire1(20, 24)    <= sub_wire18(24);
	sub_wire1(20, 25)    <= sub_wire18(25);
	sub_wire1(20, 26)    <= sub_wire18(26);
	sub_wire1(20, 27)    <= sub_wire18(27);
	sub_wire1(20, 28)    <= sub_wire18(28);
	sub_wire1(20, 29)    <= sub_wire18(29);
	sub_wire1(20, 30)    <= sub_wire18(30);
	sub_wire1(20, 31)    <= sub_wire18(31);
	sub_wire1(20, 32)    <= sub_wire18(32);
	sub_wire1(20, 33)    <= sub_wire18(33);
	sub_wire1(20, 34)    <= sub_wire18(34);
	sub_wire1(20, 35)    <= sub_wire18(35);
	sub_wire1(20, 36)    <= sub_wire18(36);
	sub_wire1(20, 37)    <= sub_wire18(37);
	sub_wire1(19, 0)    <= sub_wire19(0);
	sub_wire1(19, 1)    <= sub_wire19(1);
	sub_wire1(19, 2)    <= sub_wire19(2);
	sub_wire1(19, 3)    <= sub_wire19(3);
	sub_wire1(19, 4)    <= sub_wire19(4);
	sub_wire1(19, 5)    <= sub_wire19(5);
	sub_wire1(19, 6)    <= sub_wire19(6);
	sub_wire1(19, 7)    <= sub_wire19(7);
	sub_wire1(19, 8)    <= sub_wire19(8);
	sub_wire1(19, 9)    <= sub_wire19(9);
	sub_wire1(19, 10)    <= sub_wire19(10);
	sub_wire1(19, 11)    <= sub_wire19(11);
	sub_wire1(19, 12)    <= sub_wire19(12);
	sub_wire1(19, 13)    <= sub_wire19(13);
	sub_wire1(19, 14)    <= sub_wire19(14);
	sub_wire1(19, 15)    <= sub_wire19(15);
	sub_wire1(19, 16)    <= sub_wire19(16);
	sub_wire1(19, 17)    <= sub_wire19(17);
	sub_wire1(19, 18)    <= sub_wire19(18);
	sub_wire1(19, 19)    <= sub_wire19(19);
	sub_wire1(19, 20)    <= sub_wire19(20);
	sub_wire1(19, 21)    <= sub_wire19(21);
	sub_wire1(19, 22)    <= sub_wire19(22);
	sub_wire1(19, 23)    <= sub_wire19(23);
	sub_wire1(19, 24)    <= sub_wire19(24);
	sub_wire1(19, 25)    <= sub_wire19(25);
	sub_wire1(19, 26)    <= sub_wire19(26);
	sub_wire1(19, 27)    <= sub_wire19(27);
	sub_wire1(19, 28)    <= sub_wire19(28);
	sub_wire1(19, 29)    <= sub_wire19(29);
	sub_wire1(19, 30)    <= sub_wire19(30);
	sub_wire1(19, 31)    <= sub_wire19(31);
	sub_wire1(19, 32)    <= sub_wire19(32);
	sub_wire1(19, 33)    <= sub_wire19(33);
	sub_wire1(19, 34)    <= sub_wire19(34);
	sub_wire1(19, 35)    <= sub_wire19(35);
	sub_wire1(19, 36)    <= sub_wire19(36);
	sub_wire1(19, 37)    <= sub_wire19(37);
	sub_wire1(18, 0)    <= sub_wire20(0);
	sub_wire1(18, 1)    <= sub_wire20(1);
	sub_wire1(18, 2)    <= sub_wire20(2);
	sub_wire1(18, 3)    <= sub_wire20(3);
	sub_wire1(18, 4)    <= sub_wire20(4);
	sub_wire1(18, 5)    <= sub_wire20(5);
	sub_wire1(18, 6)    <= sub_wire20(6);
	sub_wire1(18, 7)    <= sub_wire20(7);
	sub_wire1(18, 8)    <= sub_wire20(8);
	sub_wire1(18, 9)    <= sub_wire20(9);
	sub_wire1(18, 10)    <= sub_wire20(10);
	sub_wire1(18, 11)    <= sub_wire20(11);
	sub_wire1(18, 12)    <= sub_wire20(12);
	sub_wire1(18, 13)    <= sub_wire20(13);
	sub_wire1(18, 14)    <= sub_wire20(14);
	sub_wire1(18, 15)    <= sub_wire20(15);
	sub_wire1(18, 16)    <= sub_wire20(16);
	sub_wire1(18, 17)    <= sub_wire20(17);
	sub_wire1(18, 18)    <= sub_wire20(18);
	sub_wire1(18, 19)    <= sub_wire20(19);
	sub_wire1(18, 20)    <= sub_wire20(20);
	sub_wire1(18, 21)    <= sub_wire20(21);
	sub_wire1(18, 22)    <= sub_wire20(22);
	sub_wire1(18, 23)    <= sub_wire20(23);
	sub_wire1(18, 24)    <= sub_wire20(24);
	sub_wire1(18, 25)    <= sub_wire20(25);
	sub_wire1(18, 26)    <= sub_wire20(26);
	sub_wire1(18, 27)    <= sub_wire20(27);
	sub_wire1(18, 28)    <= sub_wire20(28);
	sub_wire1(18, 29)    <= sub_wire20(29);
	sub_wire1(18, 30)    <= sub_wire20(30);
	sub_wire1(18, 31)    <= sub_wire20(31);
	sub_wire1(18, 32)    <= sub_wire20(32);
	sub_wire1(18, 33)    <= sub_wire20(33);
	sub_wire1(18, 34)    <= sub_wire20(34);
	sub_wire1(18, 35)    <= sub_wire20(35);
	sub_wire1(18, 36)    <= sub_wire20(36);
	sub_wire1(18, 37)    <= sub_wire20(37);
	sub_wire1(17, 0)    <= sub_wire21(0);
	sub_wire1(17, 1)    <= sub_wire21(1);
	sub_wire1(17, 2)    <= sub_wire21(2);
	sub_wire1(17, 3)    <= sub_wire21(3);
	sub_wire1(17, 4)    <= sub_wire21(4);
	sub_wire1(17, 5)    <= sub_wire21(5);
	sub_wire1(17, 6)    <= sub_wire21(6);
	sub_wire1(17, 7)    <= sub_wire21(7);
	sub_wire1(17, 8)    <= sub_wire21(8);
	sub_wire1(17, 9)    <= sub_wire21(9);
	sub_wire1(17, 10)    <= sub_wire21(10);
	sub_wire1(17, 11)    <= sub_wire21(11);
	sub_wire1(17, 12)    <= sub_wire21(12);
	sub_wire1(17, 13)    <= sub_wire21(13);
	sub_wire1(17, 14)    <= sub_wire21(14);
	sub_wire1(17, 15)    <= sub_wire21(15);
	sub_wire1(17, 16)    <= sub_wire21(16);
	sub_wire1(17, 17)    <= sub_wire21(17);
	sub_wire1(17, 18)    <= sub_wire21(18);
	sub_wire1(17, 19)    <= sub_wire21(19);
	sub_wire1(17, 20)    <= sub_wire21(20);
	sub_wire1(17, 21)    <= sub_wire21(21);
	sub_wire1(17, 22)    <= sub_wire21(22);
	sub_wire1(17, 23)    <= sub_wire21(23);
	sub_wire1(17, 24)    <= sub_wire21(24);
	sub_wire1(17, 25)    <= sub_wire21(25);
	sub_wire1(17, 26)    <= sub_wire21(26);
	sub_wire1(17, 27)    <= sub_wire21(27);
	sub_wire1(17, 28)    <= sub_wire21(28);
	sub_wire1(17, 29)    <= sub_wire21(29);
	sub_wire1(17, 30)    <= sub_wire21(30);
	sub_wire1(17, 31)    <= sub_wire21(31);
	sub_wire1(17, 32)    <= sub_wire21(32);
	sub_wire1(17, 33)    <= sub_wire21(33);
	sub_wire1(17, 34)    <= sub_wire21(34);
	sub_wire1(17, 35)    <= sub_wire21(35);
	sub_wire1(17, 36)    <= sub_wire21(36);
	sub_wire1(17, 37)    <= sub_wire21(37);
	sub_wire1(16, 0)    <= sub_wire22(0);
	sub_wire1(16, 1)    <= sub_wire22(1);
	sub_wire1(16, 2)    <= sub_wire22(2);
	sub_wire1(16, 3)    <= sub_wire22(3);
	sub_wire1(16, 4)    <= sub_wire22(4);
	sub_wire1(16, 5)    <= sub_wire22(5);
	sub_wire1(16, 6)    <= sub_wire22(6);
	sub_wire1(16, 7)    <= sub_wire22(7);
	sub_wire1(16, 8)    <= sub_wire22(8);
	sub_wire1(16, 9)    <= sub_wire22(9);
	sub_wire1(16, 10)    <= sub_wire22(10);
	sub_wire1(16, 11)    <= sub_wire22(11);
	sub_wire1(16, 12)    <= sub_wire22(12);
	sub_wire1(16, 13)    <= sub_wire22(13);
	sub_wire1(16, 14)    <= sub_wire22(14);
	sub_wire1(16, 15)    <= sub_wire22(15);
	sub_wire1(16, 16)    <= sub_wire22(16);
	sub_wire1(16, 17)    <= sub_wire22(17);
	sub_wire1(16, 18)    <= sub_wire22(18);
	sub_wire1(16, 19)    <= sub_wire22(19);
	sub_wire1(16, 20)    <= sub_wire22(20);
	sub_wire1(16, 21)    <= sub_wire22(21);
	sub_wire1(16, 22)    <= sub_wire22(22);
	sub_wire1(16, 23)    <= sub_wire22(23);
	sub_wire1(16, 24)    <= sub_wire22(24);
	sub_wire1(16, 25)    <= sub_wire22(25);
	sub_wire1(16, 26)    <= sub_wire22(26);
	sub_wire1(16, 27)    <= sub_wire22(27);
	sub_wire1(16, 28)    <= sub_wire22(28);
	sub_wire1(16, 29)    <= sub_wire22(29);
	sub_wire1(16, 30)    <= sub_wire22(30);
	sub_wire1(16, 31)    <= sub_wire22(31);
	sub_wire1(16, 32)    <= sub_wire22(32);
	sub_wire1(16, 33)    <= sub_wire22(33);
	sub_wire1(16, 34)    <= sub_wire22(34);
	sub_wire1(16, 35)    <= sub_wire22(35);
	sub_wire1(16, 36)    <= sub_wire22(36);
	sub_wire1(16, 37)    <= sub_wire22(37);
	sub_wire1(15, 0)    <= sub_wire23(0);
	sub_wire1(15, 1)    <= sub_wire23(1);
	sub_wire1(15, 2)    <= sub_wire23(2);
	sub_wire1(15, 3)    <= sub_wire23(3);
	sub_wire1(15, 4)    <= sub_wire23(4);
	sub_wire1(15, 5)    <= sub_wire23(5);
	sub_wire1(15, 6)    <= sub_wire23(6);
	sub_wire1(15, 7)    <= sub_wire23(7);
	sub_wire1(15, 8)    <= sub_wire23(8);
	sub_wire1(15, 9)    <= sub_wire23(9);
	sub_wire1(15, 10)    <= sub_wire23(10);
	sub_wire1(15, 11)    <= sub_wire23(11);
	sub_wire1(15, 12)    <= sub_wire23(12);
	sub_wire1(15, 13)    <= sub_wire23(13);
	sub_wire1(15, 14)    <= sub_wire23(14);
	sub_wire1(15, 15)    <= sub_wire23(15);
	sub_wire1(15, 16)    <= sub_wire23(16);
	sub_wire1(15, 17)    <= sub_wire23(17);
	sub_wire1(15, 18)    <= sub_wire23(18);
	sub_wire1(15, 19)    <= sub_wire23(19);
	sub_wire1(15, 20)    <= sub_wire23(20);
	sub_wire1(15, 21)    <= sub_wire23(21);
	sub_wire1(15, 22)    <= sub_wire23(22);
	sub_wire1(15, 23)    <= sub_wire23(23);
	sub_wire1(15, 24)    <= sub_wire23(24);
	sub_wire1(15, 25)    <= sub_wire23(25);
	sub_wire1(15, 26)    <= sub_wire23(26);
	sub_wire1(15, 27)    <= sub_wire23(27);
	sub_wire1(15, 28)    <= sub_wire23(28);
	sub_wire1(15, 29)    <= sub_wire23(29);
	sub_wire1(15, 30)    <= sub_wire23(30);
	sub_wire1(15, 31)    <= sub_wire23(31);
	sub_wire1(15, 32)    <= sub_wire23(32);
	sub_wire1(15, 33)    <= sub_wire23(33);
	sub_wire1(15, 34)    <= sub_wire23(34);
	sub_wire1(15, 35)    <= sub_wire23(35);
	sub_wire1(15, 36)    <= sub_wire23(36);
	sub_wire1(15, 37)    <= sub_wire23(37);
	sub_wire1(14, 0)    <= sub_wire24(0);
	sub_wire1(14, 1)    <= sub_wire24(1);
	sub_wire1(14, 2)    <= sub_wire24(2);
	sub_wire1(14, 3)    <= sub_wire24(3);
	sub_wire1(14, 4)    <= sub_wire24(4);
	sub_wire1(14, 5)    <= sub_wire24(5);
	sub_wire1(14, 6)    <= sub_wire24(6);
	sub_wire1(14, 7)    <= sub_wire24(7);
	sub_wire1(14, 8)    <= sub_wire24(8);
	sub_wire1(14, 9)    <= sub_wire24(9);
	sub_wire1(14, 10)    <= sub_wire24(10);
	sub_wire1(14, 11)    <= sub_wire24(11);
	sub_wire1(14, 12)    <= sub_wire24(12);
	sub_wire1(14, 13)    <= sub_wire24(13);
	sub_wire1(14, 14)    <= sub_wire24(14);
	sub_wire1(14, 15)    <= sub_wire24(15);
	sub_wire1(14, 16)    <= sub_wire24(16);
	sub_wire1(14, 17)    <= sub_wire24(17);
	sub_wire1(14, 18)    <= sub_wire24(18);
	sub_wire1(14, 19)    <= sub_wire24(19);
	sub_wire1(14, 20)    <= sub_wire24(20);
	sub_wire1(14, 21)    <= sub_wire24(21);
	sub_wire1(14, 22)    <= sub_wire24(22);
	sub_wire1(14, 23)    <= sub_wire24(23);
	sub_wire1(14, 24)    <= sub_wire24(24);
	sub_wire1(14, 25)    <= sub_wire24(25);
	sub_wire1(14, 26)    <= sub_wire24(26);
	sub_wire1(14, 27)    <= sub_wire24(27);
	sub_wire1(14, 28)    <= sub_wire24(28);
	sub_wire1(14, 29)    <= sub_wire24(29);
	sub_wire1(14, 30)    <= sub_wire24(30);
	sub_wire1(14, 31)    <= sub_wire24(31);
	sub_wire1(14, 32)    <= sub_wire24(32);
	sub_wire1(14, 33)    <= sub_wire24(33);
	sub_wire1(14, 34)    <= sub_wire24(34);
	sub_wire1(14, 35)    <= sub_wire24(35);
	sub_wire1(14, 36)    <= sub_wire24(36);
	sub_wire1(14, 37)    <= sub_wire24(37);
	sub_wire1(13, 0)    <= sub_wire25(0);
	sub_wire1(13, 1)    <= sub_wire25(1);
	sub_wire1(13, 2)    <= sub_wire25(2);
	sub_wire1(13, 3)    <= sub_wire25(3);
	sub_wire1(13, 4)    <= sub_wire25(4);
	sub_wire1(13, 5)    <= sub_wire25(5);
	sub_wire1(13, 6)    <= sub_wire25(6);
	sub_wire1(13, 7)    <= sub_wire25(7);
	sub_wire1(13, 8)    <= sub_wire25(8);
	sub_wire1(13, 9)    <= sub_wire25(9);
	sub_wire1(13, 10)    <= sub_wire25(10);
	sub_wire1(13, 11)    <= sub_wire25(11);
	sub_wire1(13, 12)    <= sub_wire25(12);
	sub_wire1(13, 13)    <= sub_wire25(13);
	sub_wire1(13, 14)    <= sub_wire25(14);
	sub_wire1(13, 15)    <= sub_wire25(15);
	sub_wire1(13, 16)    <= sub_wire25(16);
	sub_wire1(13, 17)    <= sub_wire25(17);
	sub_wire1(13, 18)    <= sub_wire25(18);
	sub_wire1(13, 19)    <= sub_wire25(19);
	sub_wire1(13, 20)    <= sub_wire25(20);
	sub_wire1(13, 21)    <= sub_wire25(21);
	sub_wire1(13, 22)    <= sub_wire25(22);
	sub_wire1(13, 23)    <= sub_wire25(23);
	sub_wire1(13, 24)    <= sub_wire25(24);
	sub_wire1(13, 25)    <= sub_wire25(25);
	sub_wire1(13, 26)    <= sub_wire25(26);
	sub_wire1(13, 27)    <= sub_wire25(27);
	sub_wire1(13, 28)    <= sub_wire25(28);
	sub_wire1(13, 29)    <= sub_wire25(29);
	sub_wire1(13, 30)    <= sub_wire25(30);
	sub_wire1(13, 31)    <= sub_wire25(31);
	sub_wire1(13, 32)    <= sub_wire25(32);
	sub_wire1(13, 33)    <= sub_wire25(33);
	sub_wire1(13, 34)    <= sub_wire25(34);
	sub_wire1(13, 35)    <= sub_wire25(35);
	sub_wire1(13, 36)    <= sub_wire25(36);
	sub_wire1(13, 37)    <= sub_wire25(37);
	sub_wire1(12, 0)    <= sub_wire26(0);
	sub_wire1(12, 1)    <= sub_wire26(1);
	sub_wire1(12, 2)    <= sub_wire26(2);
	sub_wire1(12, 3)    <= sub_wire26(3);
	sub_wire1(12, 4)    <= sub_wire26(4);
	sub_wire1(12, 5)    <= sub_wire26(5);
	sub_wire1(12, 6)    <= sub_wire26(6);
	sub_wire1(12, 7)    <= sub_wire26(7);
	sub_wire1(12, 8)    <= sub_wire26(8);
	sub_wire1(12, 9)    <= sub_wire26(9);
	sub_wire1(12, 10)    <= sub_wire26(10);
	sub_wire1(12, 11)    <= sub_wire26(11);
	sub_wire1(12, 12)    <= sub_wire26(12);
	sub_wire1(12, 13)    <= sub_wire26(13);
	sub_wire1(12, 14)    <= sub_wire26(14);
	sub_wire1(12, 15)    <= sub_wire26(15);
	sub_wire1(12, 16)    <= sub_wire26(16);
	sub_wire1(12, 17)    <= sub_wire26(17);
	sub_wire1(12, 18)    <= sub_wire26(18);
	sub_wire1(12, 19)    <= sub_wire26(19);
	sub_wire1(12, 20)    <= sub_wire26(20);
	sub_wire1(12, 21)    <= sub_wire26(21);
	sub_wire1(12, 22)    <= sub_wire26(22);
	sub_wire1(12, 23)    <= sub_wire26(23);
	sub_wire1(12, 24)    <= sub_wire26(24);
	sub_wire1(12, 25)    <= sub_wire26(25);
	sub_wire1(12, 26)    <= sub_wire26(26);
	sub_wire1(12, 27)    <= sub_wire26(27);
	sub_wire1(12, 28)    <= sub_wire26(28);
	sub_wire1(12, 29)    <= sub_wire26(29);
	sub_wire1(12, 30)    <= sub_wire26(30);
	sub_wire1(12, 31)    <= sub_wire26(31);
	sub_wire1(12, 32)    <= sub_wire26(32);
	sub_wire1(12, 33)    <= sub_wire26(33);
	sub_wire1(12, 34)    <= sub_wire26(34);
	sub_wire1(12, 35)    <= sub_wire26(35);
	sub_wire1(12, 36)    <= sub_wire26(36);
	sub_wire1(12, 37)    <= sub_wire26(37);
	sub_wire1(11, 0)    <= sub_wire27(0);
	sub_wire1(11, 1)    <= sub_wire27(1);
	sub_wire1(11, 2)    <= sub_wire27(2);
	sub_wire1(11, 3)    <= sub_wire27(3);
	sub_wire1(11, 4)    <= sub_wire27(4);
	sub_wire1(11, 5)    <= sub_wire27(5);
	sub_wire1(11, 6)    <= sub_wire27(6);
	sub_wire1(11, 7)    <= sub_wire27(7);
	sub_wire1(11, 8)    <= sub_wire27(8);
	sub_wire1(11, 9)    <= sub_wire27(9);
	sub_wire1(11, 10)    <= sub_wire27(10);
	sub_wire1(11, 11)    <= sub_wire27(11);
	sub_wire1(11, 12)    <= sub_wire27(12);
	sub_wire1(11, 13)    <= sub_wire27(13);
	sub_wire1(11, 14)    <= sub_wire27(14);
	sub_wire1(11, 15)    <= sub_wire27(15);
	sub_wire1(11, 16)    <= sub_wire27(16);
	sub_wire1(11, 17)    <= sub_wire27(17);
	sub_wire1(11, 18)    <= sub_wire27(18);
	sub_wire1(11, 19)    <= sub_wire27(19);
	sub_wire1(11, 20)    <= sub_wire27(20);
	sub_wire1(11, 21)    <= sub_wire27(21);
	sub_wire1(11, 22)    <= sub_wire27(22);
	sub_wire1(11, 23)    <= sub_wire27(23);
	sub_wire1(11, 24)    <= sub_wire27(24);
	sub_wire1(11, 25)    <= sub_wire27(25);
	sub_wire1(11, 26)    <= sub_wire27(26);
	sub_wire1(11, 27)    <= sub_wire27(27);
	sub_wire1(11, 28)    <= sub_wire27(28);
	sub_wire1(11, 29)    <= sub_wire27(29);
	sub_wire1(11, 30)    <= sub_wire27(30);
	sub_wire1(11, 31)    <= sub_wire27(31);
	sub_wire1(11, 32)    <= sub_wire27(32);
	sub_wire1(11, 33)    <= sub_wire27(33);
	sub_wire1(11, 34)    <= sub_wire27(34);
	sub_wire1(11, 35)    <= sub_wire27(35);
	sub_wire1(11, 36)    <= sub_wire27(36);
	sub_wire1(11, 37)    <= sub_wire27(37);
	sub_wire1(10, 0)    <= sub_wire28(0);
	sub_wire1(10, 1)    <= sub_wire28(1);
	sub_wire1(10, 2)    <= sub_wire28(2);
	sub_wire1(10, 3)    <= sub_wire28(3);
	sub_wire1(10, 4)    <= sub_wire28(4);
	sub_wire1(10, 5)    <= sub_wire28(5);
	sub_wire1(10, 6)    <= sub_wire28(6);
	sub_wire1(10, 7)    <= sub_wire28(7);
	sub_wire1(10, 8)    <= sub_wire28(8);
	sub_wire1(10, 9)    <= sub_wire28(9);
	sub_wire1(10, 10)    <= sub_wire28(10);
	sub_wire1(10, 11)    <= sub_wire28(11);
	sub_wire1(10, 12)    <= sub_wire28(12);
	sub_wire1(10, 13)    <= sub_wire28(13);
	sub_wire1(10, 14)    <= sub_wire28(14);
	sub_wire1(10, 15)    <= sub_wire28(15);
	sub_wire1(10, 16)    <= sub_wire28(16);
	sub_wire1(10, 17)    <= sub_wire28(17);
	sub_wire1(10, 18)    <= sub_wire28(18);
	sub_wire1(10, 19)    <= sub_wire28(19);
	sub_wire1(10, 20)    <= sub_wire28(20);
	sub_wire1(10, 21)    <= sub_wire28(21);
	sub_wire1(10, 22)    <= sub_wire28(22);
	sub_wire1(10, 23)    <= sub_wire28(23);
	sub_wire1(10, 24)    <= sub_wire28(24);
	sub_wire1(10, 25)    <= sub_wire28(25);
	sub_wire1(10, 26)    <= sub_wire28(26);
	sub_wire1(10, 27)    <= sub_wire28(27);
	sub_wire1(10, 28)    <= sub_wire28(28);
	sub_wire1(10, 29)    <= sub_wire28(29);
	sub_wire1(10, 30)    <= sub_wire28(30);
	sub_wire1(10, 31)    <= sub_wire28(31);
	sub_wire1(10, 32)    <= sub_wire28(32);
	sub_wire1(10, 33)    <= sub_wire28(33);
	sub_wire1(10, 34)    <= sub_wire28(34);
	sub_wire1(10, 35)    <= sub_wire28(35);
	sub_wire1(10, 36)    <= sub_wire28(36);
	sub_wire1(10, 37)    <= sub_wire28(37);
	sub_wire1(9, 0)    <= sub_wire29(0);
	sub_wire1(9, 1)    <= sub_wire29(1);
	sub_wire1(9, 2)    <= sub_wire29(2);
	sub_wire1(9, 3)    <= sub_wire29(3);
	sub_wire1(9, 4)    <= sub_wire29(4);
	sub_wire1(9, 5)    <= sub_wire29(5);
	sub_wire1(9, 6)    <= sub_wire29(6);
	sub_wire1(9, 7)    <= sub_wire29(7);
	sub_wire1(9, 8)    <= sub_wire29(8);
	sub_wire1(9, 9)    <= sub_wire29(9);
	sub_wire1(9, 10)    <= sub_wire29(10);
	sub_wire1(9, 11)    <= sub_wire29(11);
	sub_wire1(9, 12)    <= sub_wire29(12);
	sub_wire1(9, 13)    <= sub_wire29(13);
	sub_wire1(9, 14)    <= sub_wire29(14);
	sub_wire1(9, 15)    <= sub_wire29(15);
	sub_wire1(9, 16)    <= sub_wire29(16);
	sub_wire1(9, 17)    <= sub_wire29(17);
	sub_wire1(9, 18)    <= sub_wire29(18);
	sub_wire1(9, 19)    <= sub_wire29(19);
	sub_wire1(9, 20)    <= sub_wire29(20);
	sub_wire1(9, 21)    <= sub_wire29(21);
	sub_wire1(9, 22)    <= sub_wire29(22);
	sub_wire1(9, 23)    <= sub_wire29(23);
	sub_wire1(9, 24)    <= sub_wire29(24);
	sub_wire1(9, 25)    <= sub_wire29(25);
	sub_wire1(9, 26)    <= sub_wire29(26);
	sub_wire1(9, 27)    <= sub_wire29(27);
	sub_wire1(9, 28)    <= sub_wire29(28);
	sub_wire1(9, 29)    <= sub_wire29(29);
	sub_wire1(9, 30)    <= sub_wire29(30);
	sub_wire1(9, 31)    <= sub_wire29(31);
	sub_wire1(9, 32)    <= sub_wire29(32);
	sub_wire1(9, 33)    <= sub_wire29(33);
	sub_wire1(9, 34)    <= sub_wire29(34);
	sub_wire1(9, 35)    <= sub_wire29(35);
	sub_wire1(9, 36)    <= sub_wire29(36);
	sub_wire1(9, 37)    <= sub_wire29(37);
	sub_wire1(8, 0)    <= sub_wire30(0);
	sub_wire1(8, 1)    <= sub_wire30(1);
	sub_wire1(8, 2)    <= sub_wire30(2);
	sub_wire1(8, 3)    <= sub_wire30(3);
	sub_wire1(8, 4)    <= sub_wire30(4);
	sub_wire1(8, 5)    <= sub_wire30(5);
	sub_wire1(8, 6)    <= sub_wire30(6);
	sub_wire1(8, 7)    <= sub_wire30(7);
	sub_wire1(8, 8)    <= sub_wire30(8);
	sub_wire1(8, 9)    <= sub_wire30(9);
	sub_wire1(8, 10)    <= sub_wire30(10);
	sub_wire1(8, 11)    <= sub_wire30(11);
	sub_wire1(8, 12)    <= sub_wire30(12);
	sub_wire1(8, 13)    <= sub_wire30(13);
	sub_wire1(8, 14)    <= sub_wire30(14);
	sub_wire1(8, 15)    <= sub_wire30(15);
	sub_wire1(8, 16)    <= sub_wire30(16);
	sub_wire1(8, 17)    <= sub_wire30(17);
	sub_wire1(8, 18)    <= sub_wire30(18);
	sub_wire1(8, 19)    <= sub_wire30(19);
	sub_wire1(8, 20)    <= sub_wire30(20);
	sub_wire1(8, 21)    <= sub_wire30(21);
	sub_wire1(8, 22)    <= sub_wire30(22);
	sub_wire1(8, 23)    <= sub_wire30(23);
	sub_wire1(8, 24)    <= sub_wire30(24);
	sub_wire1(8, 25)    <= sub_wire30(25);
	sub_wire1(8, 26)    <= sub_wire30(26);
	sub_wire1(8, 27)    <= sub_wire30(27);
	sub_wire1(8, 28)    <= sub_wire30(28);
	sub_wire1(8, 29)    <= sub_wire30(29);
	sub_wire1(8, 30)    <= sub_wire30(30);
	sub_wire1(8, 31)    <= sub_wire30(31);
	sub_wire1(8, 32)    <= sub_wire30(32);
	sub_wire1(8, 33)    <= sub_wire30(33);
	sub_wire1(8, 34)    <= sub_wire30(34);
	sub_wire1(8, 35)    <= sub_wire30(35);
	sub_wire1(8, 36)    <= sub_wire30(36);
	sub_wire1(8, 37)    <= sub_wire30(37);
	sub_wire1(7, 0)    <= sub_wire31(0);
	sub_wire1(7, 1)    <= sub_wire31(1);
	sub_wire1(7, 2)    <= sub_wire31(2);
	sub_wire1(7, 3)    <= sub_wire31(3);
	sub_wire1(7, 4)    <= sub_wire31(4);
	sub_wire1(7, 5)    <= sub_wire31(5);
	sub_wire1(7, 6)    <= sub_wire31(6);
	sub_wire1(7, 7)    <= sub_wire31(7);
	sub_wire1(7, 8)    <= sub_wire31(8);
	sub_wire1(7, 9)    <= sub_wire31(9);
	sub_wire1(7, 10)    <= sub_wire31(10);
	sub_wire1(7, 11)    <= sub_wire31(11);
	sub_wire1(7, 12)    <= sub_wire31(12);
	sub_wire1(7, 13)    <= sub_wire31(13);
	sub_wire1(7, 14)    <= sub_wire31(14);
	sub_wire1(7, 15)    <= sub_wire31(15);
	sub_wire1(7, 16)    <= sub_wire31(16);
	sub_wire1(7, 17)    <= sub_wire31(17);
	sub_wire1(7, 18)    <= sub_wire31(18);
	sub_wire1(7, 19)    <= sub_wire31(19);
	sub_wire1(7, 20)    <= sub_wire31(20);
	sub_wire1(7, 21)    <= sub_wire31(21);
	sub_wire1(7, 22)    <= sub_wire31(22);
	sub_wire1(7, 23)    <= sub_wire31(23);
	sub_wire1(7, 24)    <= sub_wire31(24);
	sub_wire1(7, 25)    <= sub_wire31(25);
	sub_wire1(7, 26)    <= sub_wire31(26);
	sub_wire1(7, 27)    <= sub_wire31(27);
	sub_wire1(7, 28)    <= sub_wire31(28);
	sub_wire1(7, 29)    <= sub_wire31(29);
	sub_wire1(7, 30)    <= sub_wire31(30);
	sub_wire1(7, 31)    <= sub_wire31(31);
	sub_wire1(7, 32)    <= sub_wire31(32);
	sub_wire1(7, 33)    <= sub_wire31(33);
	sub_wire1(7, 34)    <= sub_wire31(34);
	sub_wire1(7, 35)    <= sub_wire31(35);
	sub_wire1(7, 36)    <= sub_wire31(36);
	sub_wire1(7, 37)    <= sub_wire31(37);
	sub_wire1(6, 0)    <= sub_wire32(0);
	sub_wire1(6, 1)    <= sub_wire32(1);
	sub_wire1(6, 2)    <= sub_wire32(2);
	sub_wire1(6, 3)    <= sub_wire32(3);
	sub_wire1(6, 4)    <= sub_wire32(4);
	sub_wire1(6, 5)    <= sub_wire32(5);
	sub_wire1(6, 6)    <= sub_wire32(6);
	sub_wire1(6, 7)    <= sub_wire32(7);
	sub_wire1(6, 8)    <= sub_wire32(8);
	sub_wire1(6, 9)    <= sub_wire32(9);
	sub_wire1(6, 10)    <= sub_wire32(10);
	sub_wire1(6, 11)    <= sub_wire32(11);
	sub_wire1(6, 12)    <= sub_wire32(12);
	sub_wire1(6, 13)    <= sub_wire32(13);
	sub_wire1(6, 14)    <= sub_wire32(14);
	sub_wire1(6, 15)    <= sub_wire32(15);
	sub_wire1(6, 16)    <= sub_wire32(16);
	sub_wire1(6, 17)    <= sub_wire32(17);
	sub_wire1(6, 18)    <= sub_wire32(18);
	sub_wire1(6, 19)    <= sub_wire32(19);
	sub_wire1(6, 20)    <= sub_wire32(20);
	sub_wire1(6, 21)    <= sub_wire32(21);
	sub_wire1(6, 22)    <= sub_wire32(22);
	sub_wire1(6, 23)    <= sub_wire32(23);
	sub_wire1(6, 24)    <= sub_wire32(24);
	sub_wire1(6, 25)    <= sub_wire32(25);
	sub_wire1(6, 26)    <= sub_wire32(26);
	sub_wire1(6, 27)    <= sub_wire32(27);
	sub_wire1(6, 28)    <= sub_wire32(28);
	sub_wire1(6, 29)    <= sub_wire32(29);
	sub_wire1(6, 30)    <= sub_wire32(30);
	sub_wire1(6, 31)    <= sub_wire32(31);
	sub_wire1(6, 32)    <= sub_wire32(32);
	sub_wire1(6, 33)    <= sub_wire32(33);
	sub_wire1(6, 34)    <= sub_wire32(34);
	sub_wire1(6, 35)    <= sub_wire32(35);
	sub_wire1(6, 36)    <= sub_wire32(36);
	sub_wire1(6, 37)    <= sub_wire32(37);
	sub_wire1(5, 0)    <= sub_wire33(0);
	sub_wire1(5, 1)    <= sub_wire33(1);
	sub_wire1(5, 2)    <= sub_wire33(2);
	sub_wire1(5, 3)    <= sub_wire33(3);
	sub_wire1(5, 4)    <= sub_wire33(4);
	sub_wire1(5, 5)    <= sub_wire33(5);
	sub_wire1(5, 6)    <= sub_wire33(6);
	sub_wire1(5, 7)    <= sub_wire33(7);
	sub_wire1(5, 8)    <= sub_wire33(8);
	sub_wire1(5, 9)    <= sub_wire33(9);
	sub_wire1(5, 10)    <= sub_wire33(10);
	sub_wire1(5, 11)    <= sub_wire33(11);
	sub_wire1(5, 12)    <= sub_wire33(12);
	sub_wire1(5, 13)    <= sub_wire33(13);
	sub_wire1(5, 14)    <= sub_wire33(14);
	sub_wire1(5, 15)    <= sub_wire33(15);
	sub_wire1(5, 16)    <= sub_wire33(16);
	sub_wire1(5, 17)    <= sub_wire33(17);
	sub_wire1(5, 18)    <= sub_wire33(18);
	sub_wire1(5, 19)    <= sub_wire33(19);
	sub_wire1(5, 20)    <= sub_wire33(20);
	sub_wire1(5, 21)    <= sub_wire33(21);
	sub_wire1(5, 22)    <= sub_wire33(22);
	sub_wire1(5, 23)    <= sub_wire33(23);
	sub_wire1(5, 24)    <= sub_wire33(24);
	sub_wire1(5, 25)    <= sub_wire33(25);
	sub_wire1(5, 26)    <= sub_wire33(26);
	sub_wire1(5, 27)    <= sub_wire33(27);
	sub_wire1(5, 28)    <= sub_wire33(28);
	sub_wire1(5, 29)    <= sub_wire33(29);
	sub_wire1(5, 30)    <= sub_wire33(30);
	sub_wire1(5, 31)    <= sub_wire33(31);
	sub_wire1(5, 32)    <= sub_wire33(32);
	sub_wire1(5, 33)    <= sub_wire33(33);
	sub_wire1(5, 34)    <= sub_wire33(34);
	sub_wire1(5, 35)    <= sub_wire33(35);
	sub_wire1(5, 36)    <= sub_wire33(36);
	sub_wire1(5, 37)    <= sub_wire33(37);
	sub_wire1(4, 0)    <= sub_wire34(0);
	sub_wire1(4, 1)    <= sub_wire34(1);
	sub_wire1(4, 2)    <= sub_wire34(2);
	sub_wire1(4, 3)    <= sub_wire34(3);
	sub_wire1(4, 4)    <= sub_wire34(4);
	sub_wire1(4, 5)    <= sub_wire34(5);
	sub_wire1(4, 6)    <= sub_wire34(6);
	sub_wire1(4, 7)    <= sub_wire34(7);
	sub_wire1(4, 8)    <= sub_wire34(8);
	sub_wire1(4, 9)    <= sub_wire34(9);
	sub_wire1(4, 10)    <= sub_wire34(10);
	sub_wire1(4, 11)    <= sub_wire34(11);
	sub_wire1(4, 12)    <= sub_wire34(12);
	sub_wire1(4, 13)    <= sub_wire34(13);
	sub_wire1(4, 14)    <= sub_wire34(14);
	sub_wire1(4, 15)    <= sub_wire34(15);
	sub_wire1(4, 16)    <= sub_wire34(16);
	sub_wire1(4, 17)    <= sub_wire34(17);
	sub_wire1(4, 18)    <= sub_wire34(18);
	sub_wire1(4, 19)    <= sub_wire34(19);
	sub_wire1(4, 20)    <= sub_wire34(20);
	sub_wire1(4, 21)    <= sub_wire34(21);
	sub_wire1(4, 22)    <= sub_wire34(22);
	sub_wire1(4, 23)    <= sub_wire34(23);
	sub_wire1(4, 24)    <= sub_wire34(24);
	sub_wire1(4, 25)    <= sub_wire34(25);
	sub_wire1(4, 26)    <= sub_wire34(26);
	sub_wire1(4, 27)    <= sub_wire34(27);
	sub_wire1(4, 28)    <= sub_wire34(28);
	sub_wire1(4, 29)    <= sub_wire34(29);
	sub_wire1(4, 30)    <= sub_wire34(30);
	sub_wire1(4, 31)    <= sub_wire34(31);
	sub_wire1(4, 32)    <= sub_wire34(32);
	sub_wire1(4, 33)    <= sub_wire34(33);
	sub_wire1(4, 34)    <= sub_wire34(34);
	sub_wire1(4, 35)    <= sub_wire34(35);
	sub_wire1(4, 36)    <= sub_wire34(36);
	sub_wire1(4, 37)    <= sub_wire34(37);
	sub_wire1(3, 0)    <= sub_wire35(0);
	sub_wire1(3, 1)    <= sub_wire35(1);
	sub_wire1(3, 2)    <= sub_wire35(2);
	sub_wire1(3, 3)    <= sub_wire35(3);
	sub_wire1(3, 4)    <= sub_wire35(4);
	sub_wire1(3, 5)    <= sub_wire35(5);
	sub_wire1(3, 6)    <= sub_wire35(6);
	sub_wire1(3, 7)    <= sub_wire35(7);
	sub_wire1(3, 8)    <= sub_wire35(8);
	sub_wire1(3, 9)    <= sub_wire35(9);
	sub_wire1(3, 10)    <= sub_wire35(10);
	sub_wire1(3, 11)    <= sub_wire35(11);
	sub_wire1(3, 12)    <= sub_wire35(12);
	sub_wire1(3, 13)    <= sub_wire35(13);
	sub_wire1(3, 14)    <= sub_wire35(14);
	sub_wire1(3, 15)    <= sub_wire35(15);
	sub_wire1(3, 16)    <= sub_wire35(16);
	sub_wire1(3, 17)    <= sub_wire35(17);
	sub_wire1(3, 18)    <= sub_wire35(18);
	sub_wire1(3, 19)    <= sub_wire35(19);
	sub_wire1(3, 20)    <= sub_wire35(20);
	sub_wire1(3, 21)    <= sub_wire35(21);
	sub_wire1(3, 22)    <= sub_wire35(22);
	sub_wire1(3, 23)    <= sub_wire35(23);
	sub_wire1(3, 24)    <= sub_wire35(24);
	sub_wire1(3, 25)    <= sub_wire35(25);
	sub_wire1(3, 26)    <= sub_wire35(26);
	sub_wire1(3, 27)    <= sub_wire35(27);
	sub_wire1(3, 28)    <= sub_wire35(28);
	sub_wire1(3, 29)    <= sub_wire35(29);
	sub_wire1(3, 30)    <= sub_wire35(30);
	sub_wire1(3, 31)    <= sub_wire35(31);
	sub_wire1(3, 32)    <= sub_wire35(32);
	sub_wire1(3, 33)    <= sub_wire35(33);
	sub_wire1(3, 34)    <= sub_wire35(34);
	sub_wire1(3, 35)    <= sub_wire35(35);
	sub_wire1(3, 36)    <= sub_wire35(36);
	sub_wire1(3, 37)    <= sub_wire35(37);
	sub_wire1(2, 0)    <= sub_wire36(0);
	sub_wire1(2, 1)    <= sub_wire36(1);
	sub_wire1(2, 2)    <= sub_wire36(2);
	sub_wire1(2, 3)    <= sub_wire36(3);
	sub_wire1(2, 4)    <= sub_wire36(4);
	sub_wire1(2, 5)    <= sub_wire36(5);
	sub_wire1(2, 6)    <= sub_wire36(6);
	sub_wire1(2, 7)    <= sub_wire36(7);
	sub_wire1(2, 8)    <= sub_wire36(8);
	sub_wire1(2, 9)    <= sub_wire36(9);
	sub_wire1(2, 10)    <= sub_wire36(10);
	sub_wire1(2, 11)    <= sub_wire36(11);
	sub_wire1(2, 12)    <= sub_wire36(12);
	sub_wire1(2, 13)    <= sub_wire36(13);
	sub_wire1(2, 14)    <= sub_wire36(14);
	sub_wire1(2, 15)    <= sub_wire36(15);
	sub_wire1(2, 16)    <= sub_wire36(16);
	sub_wire1(2, 17)    <= sub_wire36(17);
	sub_wire1(2, 18)    <= sub_wire36(18);
	sub_wire1(2, 19)    <= sub_wire36(19);
	sub_wire1(2, 20)    <= sub_wire36(20);
	sub_wire1(2, 21)    <= sub_wire36(21);
	sub_wire1(2, 22)    <= sub_wire36(22);
	sub_wire1(2, 23)    <= sub_wire36(23);
	sub_wire1(2, 24)    <= sub_wire36(24);
	sub_wire1(2, 25)    <= sub_wire36(25);
	sub_wire1(2, 26)    <= sub_wire36(26);
	sub_wire1(2, 27)    <= sub_wire36(27);
	sub_wire1(2, 28)    <= sub_wire36(28);
	sub_wire1(2, 29)    <= sub_wire36(29);
	sub_wire1(2, 30)    <= sub_wire36(30);
	sub_wire1(2, 31)    <= sub_wire36(31);
	sub_wire1(2, 32)    <= sub_wire36(32);
	sub_wire1(2, 33)    <= sub_wire36(33);
	sub_wire1(2, 34)    <= sub_wire36(34);
	sub_wire1(2, 35)    <= sub_wire36(35);
	sub_wire1(2, 36)    <= sub_wire36(36);
	sub_wire1(2, 37)    <= sub_wire36(37);
	sub_wire1(1, 0)    <= sub_wire37(0);
	sub_wire1(1, 1)    <= sub_wire37(1);
	sub_wire1(1, 2)    <= sub_wire37(2);
	sub_wire1(1, 3)    <= sub_wire37(3);
	sub_wire1(1, 4)    <= sub_wire37(4);
	sub_wire1(1, 5)    <= sub_wire37(5);
	sub_wire1(1, 6)    <= sub_wire37(6);
	sub_wire1(1, 7)    <= sub_wire37(7);
	sub_wire1(1, 8)    <= sub_wire37(8);
	sub_wire1(1, 9)    <= sub_wire37(9);
	sub_wire1(1, 10)    <= sub_wire37(10);
	sub_wire1(1, 11)    <= sub_wire37(11);
	sub_wire1(1, 12)    <= sub_wire37(12);
	sub_wire1(1, 13)    <= sub_wire37(13);
	sub_wire1(1, 14)    <= sub_wire37(14);
	sub_wire1(1, 15)    <= sub_wire37(15);
	sub_wire1(1, 16)    <= sub_wire37(16);
	sub_wire1(1, 17)    <= sub_wire37(17);
	sub_wire1(1, 18)    <= sub_wire37(18);
	sub_wire1(1, 19)    <= sub_wire37(19);
	sub_wire1(1, 20)    <= sub_wire37(20);
	sub_wire1(1, 21)    <= sub_wire37(21);
	sub_wire1(1, 22)    <= sub_wire37(22);
	sub_wire1(1, 23)    <= sub_wire37(23);
	sub_wire1(1, 24)    <= sub_wire37(24);
	sub_wire1(1, 25)    <= sub_wire37(25);
	sub_wire1(1, 26)    <= sub_wire37(26);
	sub_wire1(1, 27)    <= sub_wire37(27);
	sub_wire1(1, 28)    <= sub_wire37(28);
	sub_wire1(1, 29)    <= sub_wire37(29);
	sub_wire1(1, 30)    <= sub_wire37(30);
	sub_wire1(1, 31)    <= sub_wire37(31);
	sub_wire1(1, 32)    <= sub_wire37(32);
	sub_wire1(1, 33)    <= sub_wire37(33);
	sub_wire1(1, 34)    <= sub_wire37(34);
	sub_wire1(1, 35)    <= sub_wire37(35);
	sub_wire1(1, 36)    <= sub_wire37(36);
	sub_wire1(1, 37)    <= sub_wire37(37);
	sub_wire1(0, 0)    <= sub_wire38(0);
	sub_wire1(0, 1)    <= sub_wire38(1);
	sub_wire1(0, 2)    <= sub_wire38(2);
	sub_wire1(0, 3)    <= sub_wire38(3);
	sub_wire1(0, 4)    <= sub_wire38(4);
	sub_wire1(0, 5)    <= sub_wire38(5);
	sub_wire1(0, 6)    <= sub_wire38(6);
	sub_wire1(0, 7)    <= sub_wire38(7);
	sub_wire1(0, 8)    <= sub_wire38(8);
	sub_wire1(0, 9)    <= sub_wire38(9);
	sub_wire1(0, 10)    <= sub_wire38(10);
	sub_wire1(0, 11)    <= sub_wire38(11);
	sub_wire1(0, 12)    <= sub_wire38(12);
	sub_wire1(0, 13)    <= sub_wire38(13);
	sub_wire1(0, 14)    <= sub_wire38(14);
	sub_wire1(0, 15)    <= sub_wire38(15);
	sub_wire1(0, 16)    <= sub_wire38(16);
	sub_wire1(0, 17)    <= sub_wire38(17);
	sub_wire1(0, 18)    <= sub_wire38(18);
	sub_wire1(0, 19)    <= sub_wire38(19);
	sub_wire1(0, 20)    <= sub_wire38(20);
	sub_wire1(0, 21)    <= sub_wire38(21);
	sub_wire1(0, 22)    <= sub_wire38(22);
	sub_wire1(0, 23)    <= sub_wire38(23);
	sub_wire1(0, 24)    <= sub_wire38(24);
	sub_wire1(0, 25)    <= sub_wire38(25);
	sub_wire1(0, 26)    <= sub_wire38(26);
	sub_wire1(0, 27)    <= sub_wire38(27);
	sub_wire1(0, 28)    <= sub_wire38(28);
	sub_wire1(0, 29)    <= sub_wire38(29);
	sub_wire1(0, 30)    <= sub_wire38(30);
	sub_wire1(0, 31)    <= sub_wire38(31);
	sub_wire1(0, 32)    <= sub_wire38(32);
	sub_wire1(0, 33)    <= sub_wire38(33);
	sub_wire1(0, 34)    <= sub_wire38(34);
	sub_wire1(0, 35)    <= sub_wire38(35);
	sub_wire1(0, 36)    <= sub_wire38(36);
	sub_wire1(0, 37)    <= sub_wire38(37);
	result    <= sub_wire39(43 DOWNTO 0);

	parallel_add_component : parallel_add
	GENERIC MAP (
		msw_subtract => "NO",
		pipeline => 1,
		representation => "UNSIGNED",
		result_alignment => "LSB",
		shift => 0,
		size => 38,
		width => 38,
		widthr => 44,
		lpm_type => "parallel_add"
	)
	PORT MAP (
		clock => clock,
		data => sub_wire1,
		result => sub_wire39
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: MSW_SUBTRACT STRING "NO"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "1"
-- Retrieval info: CONSTANT: REPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: RESULT_ALIGNMENT STRING "LSB"
-- Retrieval info: CONSTANT: SHIFT NUMERIC "0"
-- Retrieval info: CONSTANT: SIZE NUMERIC "38"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "38"
-- Retrieval info: CONSTANT: WIDTHR NUMERIC "44"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT GND "clock"
-- Retrieval info: USED_PORT: data0x 0 0 38 0 INPUT NODEFVAL "data0x[37..0]"
-- Retrieval info: USED_PORT: data10x 0 0 38 0 INPUT NODEFVAL "data10x[37..0]"
-- Retrieval info: USED_PORT: data11x 0 0 38 0 INPUT NODEFVAL "data11x[37..0]"
-- Retrieval info: USED_PORT: data12x 0 0 38 0 INPUT NODEFVAL "data12x[37..0]"
-- Retrieval info: USED_PORT: data13x 0 0 38 0 INPUT NODEFVAL "data13x[37..0]"
-- Retrieval info: USED_PORT: data14x 0 0 38 0 INPUT NODEFVAL "data14x[37..0]"
-- Retrieval info: USED_PORT: data15x 0 0 38 0 INPUT NODEFVAL "data15x[37..0]"
-- Retrieval info: USED_PORT: data16x 0 0 38 0 INPUT NODEFVAL "data16x[37..0]"
-- Retrieval info: USED_PORT: data17x 0 0 38 0 INPUT NODEFVAL "data17x[37..0]"
-- Retrieval info: USED_PORT: data18x 0 0 38 0 INPUT NODEFVAL "data18x[37..0]"
-- Retrieval info: USED_PORT: data19x 0 0 38 0 INPUT NODEFVAL "data19x[37..0]"
-- Retrieval info: USED_PORT: data1x 0 0 38 0 INPUT NODEFVAL "data1x[37..0]"
-- Retrieval info: USED_PORT: data20x 0 0 38 0 INPUT NODEFVAL "data20x[37..0]"
-- Retrieval info: USED_PORT: data21x 0 0 38 0 INPUT NODEFVAL "data21x[37..0]"
-- Retrieval info: USED_PORT: data22x 0 0 38 0 INPUT NODEFVAL "data22x[37..0]"
-- Retrieval info: USED_PORT: data23x 0 0 38 0 INPUT NODEFVAL "data23x[37..0]"
-- Retrieval info: USED_PORT: data24x 0 0 38 0 INPUT NODEFVAL "data24x[37..0]"
-- Retrieval info: USED_PORT: data25x 0 0 38 0 INPUT NODEFVAL "data25x[37..0]"
-- Retrieval info: USED_PORT: data26x 0 0 38 0 INPUT NODEFVAL "data26x[37..0]"
-- Retrieval info: USED_PORT: data27x 0 0 38 0 INPUT NODEFVAL "data27x[37..0]"
-- Retrieval info: USED_PORT: data28x 0 0 38 0 INPUT NODEFVAL "data28x[37..0]"
-- Retrieval info: USED_PORT: data29x 0 0 38 0 INPUT NODEFVAL "data29x[37..0]"
-- Retrieval info: USED_PORT: data2x 0 0 38 0 INPUT NODEFVAL "data2x[37..0]"
-- Retrieval info: USED_PORT: data30x 0 0 38 0 INPUT NODEFVAL "data30x[37..0]"
-- Retrieval info: USED_PORT: data31x 0 0 38 0 INPUT NODEFVAL "data31x[37..0]"
-- Retrieval info: USED_PORT: data32x 0 0 38 0 INPUT NODEFVAL "data32x[37..0]"
-- Retrieval info: USED_PORT: data33x 0 0 38 0 INPUT NODEFVAL "data33x[37..0]"
-- Retrieval info: USED_PORT: data34x 0 0 38 0 INPUT NODEFVAL "data34x[37..0]"
-- Retrieval info: USED_PORT: data35x 0 0 38 0 INPUT NODEFVAL "data35x[37..0]"
-- Retrieval info: USED_PORT: data36x 0 0 38 0 INPUT NODEFVAL "data36x[37..0]"
-- Retrieval info: USED_PORT: data37x 0 0 38 0 INPUT NODEFVAL "data37x[37..0]"
-- Retrieval info: USED_PORT: data3x 0 0 38 0 INPUT NODEFVAL "data3x[37..0]"
-- Retrieval info: USED_PORT: data4x 0 0 38 0 INPUT NODEFVAL "data4x[37..0]"
-- Retrieval info: USED_PORT: data5x 0 0 38 0 INPUT NODEFVAL "data5x[37..0]"
-- Retrieval info: USED_PORT: data6x 0 0 38 0 INPUT NODEFVAL "data6x[37..0]"
-- Retrieval info: USED_PORT: data7x 0 0 38 0 INPUT NODEFVAL "data7x[37..0]"
-- Retrieval info: USED_PORT: data8x 0 0 38 0 INPUT NODEFVAL "data8x[37..0]"
-- Retrieval info: USED_PORT: data9x 0 0 38 0 INPUT NODEFVAL "data9x[37..0]"
-- Retrieval info: USED_PORT: result 0 0 44 0 OUTPUT NODEFVAL "result[43..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data 1 0 38 0 data0x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 10 38 0 data10x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 11 38 0 data11x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 12 38 0 data12x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 13 38 0 data13x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 14 38 0 data14x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 15 38 0 data15x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 16 38 0 data16x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 17 38 0 data17x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 18 38 0 data18x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 19 38 0 data19x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 1 38 0 data1x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 20 38 0 data20x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 21 38 0 data21x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 22 38 0 data22x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 23 38 0 data23x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 24 38 0 data24x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 25 38 0 data25x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 26 38 0 data26x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 27 38 0 data27x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 28 38 0 data28x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 29 38 0 data29x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 2 38 0 data2x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 30 38 0 data30x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 31 38 0 data31x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 32 38 0 data32x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 33 38 0 data33x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 34 38 0 data34x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 35 38 0 data35x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 36 38 0 data36x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 37 38 0 data37x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 3 38 0 data3x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 4 38 0 data4x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 5 38 0 data5x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 6 38 0 data6x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 7 38 0 data7x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 8 38 0 data8x 0 0 38 0
-- Retrieval info: CONNECT: @data 1 9 38 0 data9x 0 0 38 0
-- Retrieval info: CONNECT: result 0 0 44 0 @result 0 0 44 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL mapping_add.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mapping_add.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mapping_add.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mapping_add.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mapping_add_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
