-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_MUX 

-- ============================================================
-- File Name: MUX4_256b.vhd
-- Megafunction Name(s):
-- 			LPM_MUX
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 15.0.0 Build 145 04/22/2015 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus II License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY MUX4_256b IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data0x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (255 DOWNTO 0)
	);
END MUX4_256b;


ARCHITECTURE SYN OF mux4_256b IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_2D (3 DOWNTO 0, 255 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (255 DOWNTO 0);

BEGIN
	sub_wire4    <= data0x(255 DOWNTO 0);
	sub_wire3    <= data1x(255 DOWNTO 0);
	sub_wire2    <= data2x(255 DOWNTO 0);
	sub_wire0    <= data3x(255 DOWNTO 0);
	sub_wire1(3, 0)    <= sub_wire0(0);
	sub_wire1(3, 1)    <= sub_wire0(1);
	sub_wire1(3, 2)    <= sub_wire0(2);
	sub_wire1(3, 3)    <= sub_wire0(3);
	sub_wire1(3, 4)    <= sub_wire0(4);
	sub_wire1(3, 5)    <= sub_wire0(5);
	sub_wire1(3, 6)    <= sub_wire0(6);
	sub_wire1(3, 7)    <= sub_wire0(7);
	sub_wire1(3, 8)    <= sub_wire0(8);
	sub_wire1(3, 9)    <= sub_wire0(9);
	sub_wire1(3, 10)    <= sub_wire0(10);
	sub_wire1(3, 11)    <= sub_wire0(11);
	sub_wire1(3, 12)    <= sub_wire0(12);
	sub_wire1(3, 13)    <= sub_wire0(13);
	sub_wire1(3, 14)    <= sub_wire0(14);
	sub_wire1(3, 15)    <= sub_wire0(15);
	sub_wire1(3, 16)    <= sub_wire0(16);
	sub_wire1(3, 17)    <= sub_wire0(17);
	sub_wire1(3, 18)    <= sub_wire0(18);
	sub_wire1(3, 19)    <= sub_wire0(19);
	sub_wire1(3, 20)    <= sub_wire0(20);
	sub_wire1(3, 21)    <= sub_wire0(21);
	sub_wire1(3, 22)    <= sub_wire0(22);
	sub_wire1(3, 23)    <= sub_wire0(23);
	sub_wire1(3, 24)    <= sub_wire0(24);
	sub_wire1(3, 25)    <= sub_wire0(25);
	sub_wire1(3, 26)    <= sub_wire0(26);
	sub_wire1(3, 27)    <= sub_wire0(27);
	sub_wire1(3, 28)    <= sub_wire0(28);
	sub_wire1(3, 29)    <= sub_wire0(29);
	sub_wire1(3, 30)    <= sub_wire0(30);
	sub_wire1(3, 31)    <= sub_wire0(31);
	sub_wire1(3, 32)    <= sub_wire0(32);
	sub_wire1(3, 33)    <= sub_wire0(33);
	sub_wire1(3, 34)    <= sub_wire0(34);
	sub_wire1(3, 35)    <= sub_wire0(35);
	sub_wire1(3, 36)    <= sub_wire0(36);
	sub_wire1(3, 37)    <= sub_wire0(37);
	sub_wire1(3, 38)    <= sub_wire0(38);
	sub_wire1(3, 39)    <= sub_wire0(39);
	sub_wire1(3, 40)    <= sub_wire0(40);
	sub_wire1(3, 41)    <= sub_wire0(41);
	sub_wire1(3, 42)    <= sub_wire0(42);
	sub_wire1(3, 43)    <= sub_wire0(43);
	sub_wire1(3, 44)    <= sub_wire0(44);
	sub_wire1(3, 45)    <= sub_wire0(45);
	sub_wire1(3, 46)    <= sub_wire0(46);
	sub_wire1(3, 47)    <= sub_wire0(47);
	sub_wire1(3, 48)    <= sub_wire0(48);
	sub_wire1(3, 49)    <= sub_wire0(49);
	sub_wire1(3, 50)    <= sub_wire0(50);
	sub_wire1(3, 51)    <= sub_wire0(51);
	sub_wire1(3, 52)    <= sub_wire0(52);
	sub_wire1(3, 53)    <= sub_wire0(53);
	sub_wire1(3, 54)    <= sub_wire0(54);
	sub_wire1(3, 55)    <= sub_wire0(55);
	sub_wire1(3, 56)    <= sub_wire0(56);
	sub_wire1(3, 57)    <= sub_wire0(57);
	sub_wire1(3, 58)    <= sub_wire0(58);
	sub_wire1(3, 59)    <= sub_wire0(59);
	sub_wire1(3, 60)    <= sub_wire0(60);
	sub_wire1(3, 61)    <= sub_wire0(61);
	sub_wire1(3, 62)    <= sub_wire0(62);
	sub_wire1(3, 63)    <= sub_wire0(63);
	sub_wire1(3, 64)    <= sub_wire0(64);
	sub_wire1(3, 65)    <= sub_wire0(65);
	sub_wire1(3, 66)    <= sub_wire0(66);
	sub_wire1(3, 67)    <= sub_wire0(67);
	sub_wire1(3, 68)    <= sub_wire0(68);
	sub_wire1(3, 69)    <= sub_wire0(69);
	sub_wire1(3, 70)    <= sub_wire0(70);
	sub_wire1(3, 71)    <= sub_wire0(71);
	sub_wire1(3, 72)    <= sub_wire0(72);
	sub_wire1(3, 73)    <= sub_wire0(73);
	sub_wire1(3, 74)    <= sub_wire0(74);
	sub_wire1(3, 75)    <= sub_wire0(75);
	sub_wire1(3, 76)    <= sub_wire0(76);
	sub_wire1(3, 77)    <= sub_wire0(77);
	sub_wire1(3, 78)    <= sub_wire0(78);
	sub_wire1(3, 79)    <= sub_wire0(79);
	sub_wire1(3, 80)    <= sub_wire0(80);
	sub_wire1(3, 81)    <= sub_wire0(81);
	sub_wire1(3, 82)    <= sub_wire0(82);
	sub_wire1(3, 83)    <= sub_wire0(83);
	sub_wire1(3, 84)    <= sub_wire0(84);
	sub_wire1(3, 85)    <= sub_wire0(85);
	sub_wire1(3, 86)    <= sub_wire0(86);
	sub_wire1(3, 87)    <= sub_wire0(87);
	sub_wire1(3, 88)    <= sub_wire0(88);
	sub_wire1(3, 89)    <= sub_wire0(89);
	sub_wire1(3, 90)    <= sub_wire0(90);
	sub_wire1(3, 91)    <= sub_wire0(91);
	sub_wire1(3, 92)    <= sub_wire0(92);
	sub_wire1(3, 93)    <= sub_wire0(93);
	sub_wire1(3, 94)    <= sub_wire0(94);
	sub_wire1(3, 95)    <= sub_wire0(95);
	sub_wire1(3, 96)    <= sub_wire0(96);
	sub_wire1(3, 97)    <= sub_wire0(97);
	sub_wire1(3, 98)    <= sub_wire0(98);
	sub_wire1(3, 99)    <= sub_wire0(99);
	sub_wire1(3, 100)    <= sub_wire0(100);
	sub_wire1(3, 101)    <= sub_wire0(101);
	sub_wire1(3, 102)    <= sub_wire0(102);
	sub_wire1(3, 103)    <= sub_wire0(103);
	sub_wire1(3, 104)    <= sub_wire0(104);
	sub_wire1(3, 105)    <= sub_wire0(105);
	sub_wire1(3, 106)    <= sub_wire0(106);
	sub_wire1(3, 107)    <= sub_wire0(107);
	sub_wire1(3, 108)    <= sub_wire0(108);
	sub_wire1(3, 109)    <= sub_wire0(109);
	sub_wire1(3, 110)    <= sub_wire0(110);
	sub_wire1(3, 111)    <= sub_wire0(111);
	sub_wire1(3, 112)    <= sub_wire0(112);
	sub_wire1(3, 113)    <= sub_wire0(113);
	sub_wire1(3, 114)    <= sub_wire0(114);
	sub_wire1(3, 115)    <= sub_wire0(115);
	sub_wire1(3, 116)    <= sub_wire0(116);
	sub_wire1(3, 117)    <= sub_wire0(117);
	sub_wire1(3, 118)    <= sub_wire0(118);
	sub_wire1(3, 119)    <= sub_wire0(119);
	sub_wire1(3, 120)    <= sub_wire0(120);
	sub_wire1(3, 121)    <= sub_wire0(121);
	sub_wire1(3, 122)    <= sub_wire0(122);
	sub_wire1(3, 123)    <= sub_wire0(123);
	sub_wire1(3, 124)    <= sub_wire0(124);
	sub_wire1(3, 125)    <= sub_wire0(125);
	sub_wire1(3, 126)    <= sub_wire0(126);
	sub_wire1(3, 127)    <= sub_wire0(127);
	sub_wire1(3, 128)    <= sub_wire0(128);
	sub_wire1(3, 129)    <= sub_wire0(129);
	sub_wire1(3, 130)    <= sub_wire0(130);
	sub_wire1(3, 131)    <= sub_wire0(131);
	sub_wire1(3, 132)    <= sub_wire0(132);
	sub_wire1(3, 133)    <= sub_wire0(133);
	sub_wire1(3, 134)    <= sub_wire0(134);
	sub_wire1(3, 135)    <= sub_wire0(135);
	sub_wire1(3, 136)    <= sub_wire0(136);
	sub_wire1(3, 137)    <= sub_wire0(137);
	sub_wire1(3, 138)    <= sub_wire0(138);
	sub_wire1(3, 139)    <= sub_wire0(139);
	sub_wire1(3, 140)    <= sub_wire0(140);
	sub_wire1(3, 141)    <= sub_wire0(141);
	sub_wire1(3, 142)    <= sub_wire0(142);
	sub_wire1(3, 143)    <= sub_wire0(143);
	sub_wire1(3, 144)    <= sub_wire0(144);
	sub_wire1(3, 145)    <= sub_wire0(145);
	sub_wire1(3, 146)    <= sub_wire0(146);
	sub_wire1(3, 147)    <= sub_wire0(147);
	sub_wire1(3, 148)    <= sub_wire0(148);
	sub_wire1(3, 149)    <= sub_wire0(149);
	sub_wire1(3, 150)    <= sub_wire0(150);
	sub_wire1(3, 151)    <= sub_wire0(151);
	sub_wire1(3, 152)    <= sub_wire0(152);
	sub_wire1(3, 153)    <= sub_wire0(153);
	sub_wire1(3, 154)    <= sub_wire0(154);
	sub_wire1(3, 155)    <= sub_wire0(155);
	sub_wire1(3, 156)    <= sub_wire0(156);
	sub_wire1(3, 157)    <= sub_wire0(157);
	sub_wire1(3, 158)    <= sub_wire0(158);
	sub_wire1(3, 159)    <= sub_wire0(159);
	sub_wire1(3, 160)    <= sub_wire0(160);
	sub_wire1(3, 161)    <= sub_wire0(161);
	sub_wire1(3, 162)    <= sub_wire0(162);
	sub_wire1(3, 163)    <= sub_wire0(163);
	sub_wire1(3, 164)    <= sub_wire0(164);
	sub_wire1(3, 165)    <= sub_wire0(165);
	sub_wire1(3, 166)    <= sub_wire0(166);
	sub_wire1(3, 167)    <= sub_wire0(167);
	sub_wire1(3, 168)    <= sub_wire0(168);
	sub_wire1(3, 169)    <= sub_wire0(169);
	sub_wire1(3, 170)    <= sub_wire0(170);
	sub_wire1(3, 171)    <= sub_wire0(171);
	sub_wire1(3, 172)    <= sub_wire0(172);
	sub_wire1(3, 173)    <= sub_wire0(173);
	sub_wire1(3, 174)    <= sub_wire0(174);
	sub_wire1(3, 175)    <= sub_wire0(175);
	sub_wire1(3, 176)    <= sub_wire0(176);
	sub_wire1(3, 177)    <= sub_wire0(177);
	sub_wire1(3, 178)    <= sub_wire0(178);
	sub_wire1(3, 179)    <= sub_wire0(179);
	sub_wire1(3, 180)    <= sub_wire0(180);
	sub_wire1(3, 181)    <= sub_wire0(181);
	sub_wire1(3, 182)    <= sub_wire0(182);
	sub_wire1(3, 183)    <= sub_wire0(183);
	sub_wire1(3, 184)    <= sub_wire0(184);
	sub_wire1(3, 185)    <= sub_wire0(185);
	sub_wire1(3, 186)    <= sub_wire0(186);
	sub_wire1(3, 187)    <= sub_wire0(187);
	sub_wire1(3, 188)    <= sub_wire0(188);
	sub_wire1(3, 189)    <= sub_wire0(189);
	sub_wire1(3, 190)    <= sub_wire0(190);
	sub_wire1(3, 191)    <= sub_wire0(191);
	sub_wire1(3, 192)    <= sub_wire0(192);
	sub_wire1(3, 193)    <= sub_wire0(193);
	sub_wire1(3, 194)    <= sub_wire0(194);
	sub_wire1(3, 195)    <= sub_wire0(195);
	sub_wire1(3, 196)    <= sub_wire0(196);
	sub_wire1(3, 197)    <= sub_wire0(197);
	sub_wire1(3, 198)    <= sub_wire0(198);
	sub_wire1(3, 199)    <= sub_wire0(199);
	sub_wire1(3, 200)    <= sub_wire0(200);
	sub_wire1(3, 201)    <= sub_wire0(201);
	sub_wire1(3, 202)    <= sub_wire0(202);
	sub_wire1(3, 203)    <= sub_wire0(203);
	sub_wire1(3, 204)    <= sub_wire0(204);
	sub_wire1(3, 205)    <= sub_wire0(205);
	sub_wire1(3, 206)    <= sub_wire0(206);
	sub_wire1(3, 207)    <= sub_wire0(207);
	sub_wire1(3, 208)    <= sub_wire0(208);
	sub_wire1(3, 209)    <= sub_wire0(209);
	sub_wire1(3, 210)    <= sub_wire0(210);
	sub_wire1(3, 211)    <= sub_wire0(211);
	sub_wire1(3, 212)    <= sub_wire0(212);
	sub_wire1(3, 213)    <= sub_wire0(213);
	sub_wire1(3, 214)    <= sub_wire0(214);
	sub_wire1(3, 215)    <= sub_wire0(215);
	sub_wire1(3, 216)    <= sub_wire0(216);
	sub_wire1(3, 217)    <= sub_wire0(217);
	sub_wire1(3, 218)    <= sub_wire0(218);
	sub_wire1(3, 219)    <= sub_wire0(219);
	sub_wire1(3, 220)    <= sub_wire0(220);
	sub_wire1(3, 221)    <= sub_wire0(221);
	sub_wire1(3, 222)    <= sub_wire0(222);
	sub_wire1(3, 223)    <= sub_wire0(223);
	sub_wire1(3, 224)    <= sub_wire0(224);
	sub_wire1(3, 225)    <= sub_wire0(225);
	sub_wire1(3, 226)    <= sub_wire0(226);
	sub_wire1(3, 227)    <= sub_wire0(227);
	sub_wire1(3, 228)    <= sub_wire0(228);
	sub_wire1(3, 229)    <= sub_wire0(229);
	sub_wire1(3, 230)    <= sub_wire0(230);
	sub_wire1(3, 231)    <= sub_wire0(231);
	sub_wire1(3, 232)    <= sub_wire0(232);
	sub_wire1(3, 233)    <= sub_wire0(233);
	sub_wire1(3, 234)    <= sub_wire0(234);
	sub_wire1(3, 235)    <= sub_wire0(235);
	sub_wire1(3, 236)    <= sub_wire0(236);
	sub_wire1(3, 237)    <= sub_wire0(237);
	sub_wire1(3, 238)    <= sub_wire0(238);
	sub_wire1(3, 239)    <= sub_wire0(239);
	sub_wire1(3, 240)    <= sub_wire0(240);
	sub_wire1(3, 241)    <= sub_wire0(241);
	sub_wire1(3, 242)    <= sub_wire0(242);
	sub_wire1(3, 243)    <= sub_wire0(243);
	sub_wire1(3, 244)    <= sub_wire0(244);
	sub_wire1(3, 245)    <= sub_wire0(245);
	sub_wire1(3, 246)    <= sub_wire0(246);
	sub_wire1(3, 247)    <= sub_wire0(247);
	sub_wire1(3, 248)    <= sub_wire0(248);
	sub_wire1(3, 249)    <= sub_wire0(249);
	sub_wire1(3, 250)    <= sub_wire0(250);
	sub_wire1(3, 251)    <= sub_wire0(251);
	sub_wire1(3, 252)    <= sub_wire0(252);
	sub_wire1(3, 253)    <= sub_wire0(253);
	sub_wire1(3, 254)    <= sub_wire0(254);
	sub_wire1(3, 255)    <= sub_wire0(255);
	sub_wire1(2, 0)    <= sub_wire2(0);
	sub_wire1(2, 1)    <= sub_wire2(1);
	sub_wire1(2, 2)    <= sub_wire2(2);
	sub_wire1(2, 3)    <= sub_wire2(3);
	sub_wire1(2, 4)    <= sub_wire2(4);
	sub_wire1(2, 5)    <= sub_wire2(5);
	sub_wire1(2, 6)    <= sub_wire2(6);
	sub_wire1(2, 7)    <= sub_wire2(7);
	sub_wire1(2, 8)    <= sub_wire2(8);
	sub_wire1(2, 9)    <= sub_wire2(9);
	sub_wire1(2, 10)    <= sub_wire2(10);
	sub_wire1(2, 11)    <= sub_wire2(11);
	sub_wire1(2, 12)    <= sub_wire2(12);
	sub_wire1(2, 13)    <= sub_wire2(13);
	sub_wire1(2, 14)    <= sub_wire2(14);
	sub_wire1(2, 15)    <= sub_wire2(15);
	sub_wire1(2, 16)    <= sub_wire2(16);
	sub_wire1(2, 17)    <= sub_wire2(17);
	sub_wire1(2, 18)    <= sub_wire2(18);
	sub_wire1(2, 19)    <= sub_wire2(19);
	sub_wire1(2, 20)    <= sub_wire2(20);
	sub_wire1(2, 21)    <= sub_wire2(21);
	sub_wire1(2, 22)    <= sub_wire2(22);
	sub_wire1(2, 23)    <= sub_wire2(23);
	sub_wire1(2, 24)    <= sub_wire2(24);
	sub_wire1(2, 25)    <= sub_wire2(25);
	sub_wire1(2, 26)    <= sub_wire2(26);
	sub_wire1(2, 27)    <= sub_wire2(27);
	sub_wire1(2, 28)    <= sub_wire2(28);
	sub_wire1(2, 29)    <= sub_wire2(29);
	sub_wire1(2, 30)    <= sub_wire2(30);
	sub_wire1(2, 31)    <= sub_wire2(31);
	sub_wire1(2, 32)    <= sub_wire2(32);
	sub_wire1(2, 33)    <= sub_wire2(33);
	sub_wire1(2, 34)    <= sub_wire2(34);
	sub_wire1(2, 35)    <= sub_wire2(35);
	sub_wire1(2, 36)    <= sub_wire2(36);
	sub_wire1(2, 37)    <= sub_wire2(37);
	sub_wire1(2, 38)    <= sub_wire2(38);
	sub_wire1(2, 39)    <= sub_wire2(39);
	sub_wire1(2, 40)    <= sub_wire2(40);
	sub_wire1(2, 41)    <= sub_wire2(41);
	sub_wire1(2, 42)    <= sub_wire2(42);
	sub_wire1(2, 43)    <= sub_wire2(43);
	sub_wire1(2, 44)    <= sub_wire2(44);
	sub_wire1(2, 45)    <= sub_wire2(45);
	sub_wire1(2, 46)    <= sub_wire2(46);
	sub_wire1(2, 47)    <= sub_wire2(47);
	sub_wire1(2, 48)    <= sub_wire2(48);
	sub_wire1(2, 49)    <= sub_wire2(49);
	sub_wire1(2, 50)    <= sub_wire2(50);
	sub_wire1(2, 51)    <= sub_wire2(51);
	sub_wire1(2, 52)    <= sub_wire2(52);
	sub_wire1(2, 53)    <= sub_wire2(53);
	sub_wire1(2, 54)    <= sub_wire2(54);
	sub_wire1(2, 55)    <= sub_wire2(55);
	sub_wire1(2, 56)    <= sub_wire2(56);
	sub_wire1(2, 57)    <= sub_wire2(57);
	sub_wire1(2, 58)    <= sub_wire2(58);
	sub_wire1(2, 59)    <= sub_wire2(59);
	sub_wire1(2, 60)    <= sub_wire2(60);
	sub_wire1(2, 61)    <= sub_wire2(61);
	sub_wire1(2, 62)    <= sub_wire2(62);
	sub_wire1(2, 63)    <= sub_wire2(63);
	sub_wire1(2, 64)    <= sub_wire2(64);
	sub_wire1(2, 65)    <= sub_wire2(65);
	sub_wire1(2, 66)    <= sub_wire2(66);
	sub_wire1(2, 67)    <= sub_wire2(67);
	sub_wire1(2, 68)    <= sub_wire2(68);
	sub_wire1(2, 69)    <= sub_wire2(69);
	sub_wire1(2, 70)    <= sub_wire2(70);
	sub_wire1(2, 71)    <= sub_wire2(71);
	sub_wire1(2, 72)    <= sub_wire2(72);
	sub_wire1(2, 73)    <= sub_wire2(73);
	sub_wire1(2, 74)    <= sub_wire2(74);
	sub_wire1(2, 75)    <= sub_wire2(75);
	sub_wire1(2, 76)    <= sub_wire2(76);
	sub_wire1(2, 77)    <= sub_wire2(77);
	sub_wire1(2, 78)    <= sub_wire2(78);
	sub_wire1(2, 79)    <= sub_wire2(79);
	sub_wire1(2, 80)    <= sub_wire2(80);
	sub_wire1(2, 81)    <= sub_wire2(81);
	sub_wire1(2, 82)    <= sub_wire2(82);
	sub_wire1(2, 83)    <= sub_wire2(83);
	sub_wire1(2, 84)    <= sub_wire2(84);
	sub_wire1(2, 85)    <= sub_wire2(85);
	sub_wire1(2, 86)    <= sub_wire2(86);
	sub_wire1(2, 87)    <= sub_wire2(87);
	sub_wire1(2, 88)    <= sub_wire2(88);
	sub_wire1(2, 89)    <= sub_wire2(89);
	sub_wire1(2, 90)    <= sub_wire2(90);
	sub_wire1(2, 91)    <= sub_wire2(91);
	sub_wire1(2, 92)    <= sub_wire2(92);
	sub_wire1(2, 93)    <= sub_wire2(93);
	sub_wire1(2, 94)    <= sub_wire2(94);
	sub_wire1(2, 95)    <= sub_wire2(95);
	sub_wire1(2, 96)    <= sub_wire2(96);
	sub_wire1(2, 97)    <= sub_wire2(97);
	sub_wire1(2, 98)    <= sub_wire2(98);
	sub_wire1(2, 99)    <= sub_wire2(99);
	sub_wire1(2, 100)    <= sub_wire2(100);
	sub_wire1(2, 101)    <= sub_wire2(101);
	sub_wire1(2, 102)    <= sub_wire2(102);
	sub_wire1(2, 103)    <= sub_wire2(103);
	sub_wire1(2, 104)    <= sub_wire2(104);
	sub_wire1(2, 105)    <= sub_wire2(105);
	sub_wire1(2, 106)    <= sub_wire2(106);
	sub_wire1(2, 107)    <= sub_wire2(107);
	sub_wire1(2, 108)    <= sub_wire2(108);
	sub_wire1(2, 109)    <= sub_wire2(109);
	sub_wire1(2, 110)    <= sub_wire2(110);
	sub_wire1(2, 111)    <= sub_wire2(111);
	sub_wire1(2, 112)    <= sub_wire2(112);
	sub_wire1(2, 113)    <= sub_wire2(113);
	sub_wire1(2, 114)    <= sub_wire2(114);
	sub_wire1(2, 115)    <= sub_wire2(115);
	sub_wire1(2, 116)    <= sub_wire2(116);
	sub_wire1(2, 117)    <= sub_wire2(117);
	sub_wire1(2, 118)    <= sub_wire2(118);
	sub_wire1(2, 119)    <= sub_wire2(119);
	sub_wire1(2, 120)    <= sub_wire2(120);
	sub_wire1(2, 121)    <= sub_wire2(121);
	sub_wire1(2, 122)    <= sub_wire2(122);
	sub_wire1(2, 123)    <= sub_wire2(123);
	sub_wire1(2, 124)    <= sub_wire2(124);
	sub_wire1(2, 125)    <= sub_wire2(125);
	sub_wire1(2, 126)    <= sub_wire2(126);
	sub_wire1(2, 127)    <= sub_wire2(127);
	sub_wire1(2, 128)    <= sub_wire2(128);
	sub_wire1(2, 129)    <= sub_wire2(129);
	sub_wire1(2, 130)    <= sub_wire2(130);
	sub_wire1(2, 131)    <= sub_wire2(131);
	sub_wire1(2, 132)    <= sub_wire2(132);
	sub_wire1(2, 133)    <= sub_wire2(133);
	sub_wire1(2, 134)    <= sub_wire2(134);
	sub_wire1(2, 135)    <= sub_wire2(135);
	sub_wire1(2, 136)    <= sub_wire2(136);
	sub_wire1(2, 137)    <= sub_wire2(137);
	sub_wire1(2, 138)    <= sub_wire2(138);
	sub_wire1(2, 139)    <= sub_wire2(139);
	sub_wire1(2, 140)    <= sub_wire2(140);
	sub_wire1(2, 141)    <= sub_wire2(141);
	sub_wire1(2, 142)    <= sub_wire2(142);
	sub_wire1(2, 143)    <= sub_wire2(143);
	sub_wire1(2, 144)    <= sub_wire2(144);
	sub_wire1(2, 145)    <= sub_wire2(145);
	sub_wire1(2, 146)    <= sub_wire2(146);
	sub_wire1(2, 147)    <= sub_wire2(147);
	sub_wire1(2, 148)    <= sub_wire2(148);
	sub_wire1(2, 149)    <= sub_wire2(149);
	sub_wire1(2, 150)    <= sub_wire2(150);
	sub_wire1(2, 151)    <= sub_wire2(151);
	sub_wire1(2, 152)    <= sub_wire2(152);
	sub_wire1(2, 153)    <= sub_wire2(153);
	sub_wire1(2, 154)    <= sub_wire2(154);
	sub_wire1(2, 155)    <= sub_wire2(155);
	sub_wire1(2, 156)    <= sub_wire2(156);
	sub_wire1(2, 157)    <= sub_wire2(157);
	sub_wire1(2, 158)    <= sub_wire2(158);
	sub_wire1(2, 159)    <= sub_wire2(159);
	sub_wire1(2, 160)    <= sub_wire2(160);
	sub_wire1(2, 161)    <= sub_wire2(161);
	sub_wire1(2, 162)    <= sub_wire2(162);
	sub_wire1(2, 163)    <= sub_wire2(163);
	sub_wire1(2, 164)    <= sub_wire2(164);
	sub_wire1(2, 165)    <= sub_wire2(165);
	sub_wire1(2, 166)    <= sub_wire2(166);
	sub_wire1(2, 167)    <= sub_wire2(167);
	sub_wire1(2, 168)    <= sub_wire2(168);
	sub_wire1(2, 169)    <= sub_wire2(169);
	sub_wire1(2, 170)    <= sub_wire2(170);
	sub_wire1(2, 171)    <= sub_wire2(171);
	sub_wire1(2, 172)    <= sub_wire2(172);
	sub_wire1(2, 173)    <= sub_wire2(173);
	sub_wire1(2, 174)    <= sub_wire2(174);
	sub_wire1(2, 175)    <= sub_wire2(175);
	sub_wire1(2, 176)    <= sub_wire2(176);
	sub_wire1(2, 177)    <= sub_wire2(177);
	sub_wire1(2, 178)    <= sub_wire2(178);
	sub_wire1(2, 179)    <= sub_wire2(179);
	sub_wire1(2, 180)    <= sub_wire2(180);
	sub_wire1(2, 181)    <= sub_wire2(181);
	sub_wire1(2, 182)    <= sub_wire2(182);
	sub_wire1(2, 183)    <= sub_wire2(183);
	sub_wire1(2, 184)    <= sub_wire2(184);
	sub_wire1(2, 185)    <= sub_wire2(185);
	sub_wire1(2, 186)    <= sub_wire2(186);
	sub_wire1(2, 187)    <= sub_wire2(187);
	sub_wire1(2, 188)    <= sub_wire2(188);
	sub_wire1(2, 189)    <= sub_wire2(189);
	sub_wire1(2, 190)    <= sub_wire2(190);
	sub_wire1(2, 191)    <= sub_wire2(191);
	sub_wire1(2, 192)    <= sub_wire2(192);
	sub_wire1(2, 193)    <= sub_wire2(193);
	sub_wire1(2, 194)    <= sub_wire2(194);
	sub_wire1(2, 195)    <= sub_wire2(195);
	sub_wire1(2, 196)    <= sub_wire2(196);
	sub_wire1(2, 197)    <= sub_wire2(197);
	sub_wire1(2, 198)    <= sub_wire2(198);
	sub_wire1(2, 199)    <= sub_wire2(199);
	sub_wire1(2, 200)    <= sub_wire2(200);
	sub_wire1(2, 201)    <= sub_wire2(201);
	sub_wire1(2, 202)    <= sub_wire2(202);
	sub_wire1(2, 203)    <= sub_wire2(203);
	sub_wire1(2, 204)    <= sub_wire2(204);
	sub_wire1(2, 205)    <= sub_wire2(205);
	sub_wire1(2, 206)    <= sub_wire2(206);
	sub_wire1(2, 207)    <= sub_wire2(207);
	sub_wire1(2, 208)    <= sub_wire2(208);
	sub_wire1(2, 209)    <= sub_wire2(209);
	sub_wire1(2, 210)    <= sub_wire2(210);
	sub_wire1(2, 211)    <= sub_wire2(211);
	sub_wire1(2, 212)    <= sub_wire2(212);
	sub_wire1(2, 213)    <= sub_wire2(213);
	sub_wire1(2, 214)    <= sub_wire2(214);
	sub_wire1(2, 215)    <= sub_wire2(215);
	sub_wire1(2, 216)    <= sub_wire2(216);
	sub_wire1(2, 217)    <= sub_wire2(217);
	sub_wire1(2, 218)    <= sub_wire2(218);
	sub_wire1(2, 219)    <= sub_wire2(219);
	sub_wire1(2, 220)    <= sub_wire2(220);
	sub_wire1(2, 221)    <= sub_wire2(221);
	sub_wire1(2, 222)    <= sub_wire2(222);
	sub_wire1(2, 223)    <= sub_wire2(223);
	sub_wire1(2, 224)    <= sub_wire2(224);
	sub_wire1(2, 225)    <= sub_wire2(225);
	sub_wire1(2, 226)    <= sub_wire2(226);
	sub_wire1(2, 227)    <= sub_wire2(227);
	sub_wire1(2, 228)    <= sub_wire2(228);
	sub_wire1(2, 229)    <= sub_wire2(229);
	sub_wire1(2, 230)    <= sub_wire2(230);
	sub_wire1(2, 231)    <= sub_wire2(231);
	sub_wire1(2, 232)    <= sub_wire2(232);
	sub_wire1(2, 233)    <= sub_wire2(233);
	sub_wire1(2, 234)    <= sub_wire2(234);
	sub_wire1(2, 235)    <= sub_wire2(235);
	sub_wire1(2, 236)    <= sub_wire2(236);
	sub_wire1(2, 237)    <= sub_wire2(237);
	sub_wire1(2, 238)    <= sub_wire2(238);
	sub_wire1(2, 239)    <= sub_wire2(239);
	sub_wire1(2, 240)    <= sub_wire2(240);
	sub_wire1(2, 241)    <= sub_wire2(241);
	sub_wire1(2, 242)    <= sub_wire2(242);
	sub_wire1(2, 243)    <= sub_wire2(243);
	sub_wire1(2, 244)    <= sub_wire2(244);
	sub_wire1(2, 245)    <= sub_wire2(245);
	sub_wire1(2, 246)    <= sub_wire2(246);
	sub_wire1(2, 247)    <= sub_wire2(247);
	sub_wire1(2, 248)    <= sub_wire2(248);
	sub_wire1(2, 249)    <= sub_wire2(249);
	sub_wire1(2, 250)    <= sub_wire2(250);
	sub_wire1(2, 251)    <= sub_wire2(251);
	sub_wire1(2, 252)    <= sub_wire2(252);
	sub_wire1(2, 253)    <= sub_wire2(253);
	sub_wire1(2, 254)    <= sub_wire2(254);
	sub_wire1(2, 255)    <= sub_wire2(255);
	sub_wire1(1, 0)    <= sub_wire3(0);
	sub_wire1(1, 1)    <= sub_wire3(1);
	sub_wire1(1, 2)    <= sub_wire3(2);
	sub_wire1(1, 3)    <= sub_wire3(3);
	sub_wire1(1, 4)    <= sub_wire3(4);
	sub_wire1(1, 5)    <= sub_wire3(5);
	sub_wire1(1, 6)    <= sub_wire3(6);
	sub_wire1(1, 7)    <= sub_wire3(7);
	sub_wire1(1, 8)    <= sub_wire3(8);
	sub_wire1(1, 9)    <= sub_wire3(9);
	sub_wire1(1, 10)    <= sub_wire3(10);
	sub_wire1(1, 11)    <= sub_wire3(11);
	sub_wire1(1, 12)    <= sub_wire3(12);
	sub_wire1(1, 13)    <= sub_wire3(13);
	sub_wire1(1, 14)    <= sub_wire3(14);
	sub_wire1(1, 15)    <= sub_wire3(15);
	sub_wire1(1, 16)    <= sub_wire3(16);
	sub_wire1(1, 17)    <= sub_wire3(17);
	sub_wire1(1, 18)    <= sub_wire3(18);
	sub_wire1(1, 19)    <= sub_wire3(19);
	sub_wire1(1, 20)    <= sub_wire3(20);
	sub_wire1(1, 21)    <= sub_wire3(21);
	sub_wire1(1, 22)    <= sub_wire3(22);
	sub_wire1(1, 23)    <= sub_wire3(23);
	sub_wire1(1, 24)    <= sub_wire3(24);
	sub_wire1(1, 25)    <= sub_wire3(25);
	sub_wire1(1, 26)    <= sub_wire3(26);
	sub_wire1(1, 27)    <= sub_wire3(27);
	sub_wire1(1, 28)    <= sub_wire3(28);
	sub_wire1(1, 29)    <= sub_wire3(29);
	sub_wire1(1, 30)    <= sub_wire3(30);
	sub_wire1(1, 31)    <= sub_wire3(31);
	sub_wire1(1, 32)    <= sub_wire3(32);
	sub_wire1(1, 33)    <= sub_wire3(33);
	sub_wire1(1, 34)    <= sub_wire3(34);
	sub_wire1(1, 35)    <= sub_wire3(35);
	sub_wire1(1, 36)    <= sub_wire3(36);
	sub_wire1(1, 37)    <= sub_wire3(37);
	sub_wire1(1, 38)    <= sub_wire3(38);
	sub_wire1(1, 39)    <= sub_wire3(39);
	sub_wire1(1, 40)    <= sub_wire3(40);
	sub_wire1(1, 41)    <= sub_wire3(41);
	sub_wire1(1, 42)    <= sub_wire3(42);
	sub_wire1(1, 43)    <= sub_wire3(43);
	sub_wire1(1, 44)    <= sub_wire3(44);
	sub_wire1(1, 45)    <= sub_wire3(45);
	sub_wire1(1, 46)    <= sub_wire3(46);
	sub_wire1(1, 47)    <= sub_wire3(47);
	sub_wire1(1, 48)    <= sub_wire3(48);
	sub_wire1(1, 49)    <= sub_wire3(49);
	sub_wire1(1, 50)    <= sub_wire3(50);
	sub_wire1(1, 51)    <= sub_wire3(51);
	sub_wire1(1, 52)    <= sub_wire3(52);
	sub_wire1(1, 53)    <= sub_wire3(53);
	sub_wire1(1, 54)    <= sub_wire3(54);
	sub_wire1(1, 55)    <= sub_wire3(55);
	sub_wire1(1, 56)    <= sub_wire3(56);
	sub_wire1(1, 57)    <= sub_wire3(57);
	sub_wire1(1, 58)    <= sub_wire3(58);
	sub_wire1(1, 59)    <= sub_wire3(59);
	sub_wire1(1, 60)    <= sub_wire3(60);
	sub_wire1(1, 61)    <= sub_wire3(61);
	sub_wire1(1, 62)    <= sub_wire3(62);
	sub_wire1(1, 63)    <= sub_wire3(63);
	sub_wire1(1, 64)    <= sub_wire3(64);
	sub_wire1(1, 65)    <= sub_wire3(65);
	sub_wire1(1, 66)    <= sub_wire3(66);
	sub_wire1(1, 67)    <= sub_wire3(67);
	sub_wire1(1, 68)    <= sub_wire3(68);
	sub_wire1(1, 69)    <= sub_wire3(69);
	sub_wire1(1, 70)    <= sub_wire3(70);
	sub_wire1(1, 71)    <= sub_wire3(71);
	sub_wire1(1, 72)    <= sub_wire3(72);
	sub_wire1(1, 73)    <= sub_wire3(73);
	sub_wire1(1, 74)    <= sub_wire3(74);
	sub_wire1(1, 75)    <= sub_wire3(75);
	sub_wire1(1, 76)    <= sub_wire3(76);
	sub_wire1(1, 77)    <= sub_wire3(77);
	sub_wire1(1, 78)    <= sub_wire3(78);
	sub_wire1(1, 79)    <= sub_wire3(79);
	sub_wire1(1, 80)    <= sub_wire3(80);
	sub_wire1(1, 81)    <= sub_wire3(81);
	sub_wire1(1, 82)    <= sub_wire3(82);
	sub_wire1(1, 83)    <= sub_wire3(83);
	sub_wire1(1, 84)    <= sub_wire3(84);
	sub_wire1(1, 85)    <= sub_wire3(85);
	sub_wire1(1, 86)    <= sub_wire3(86);
	sub_wire1(1, 87)    <= sub_wire3(87);
	sub_wire1(1, 88)    <= sub_wire3(88);
	sub_wire1(1, 89)    <= sub_wire3(89);
	sub_wire1(1, 90)    <= sub_wire3(90);
	sub_wire1(1, 91)    <= sub_wire3(91);
	sub_wire1(1, 92)    <= sub_wire3(92);
	sub_wire1(1, 93)    <= sub_wire3(93);
	sub_wire1(1, 94)    <= sub_wire3(94);
	sub_wire1(1, 95)    <= sub_wire3(95);
	sub_wire1(1, 96)    <= sub_wire3(96);
	sub_wire1(1, 97)    <= sub_wire3(97);
	sub_wire1(1, 98)    <= sub_wire3(98);
	sub_wire1(1, 99)    <= sub_wire3(99);
	sub_wire1(1, 100)    <= sub_wire3(100);
	sub_wire1(1, 101)    <= sub_wire3(101);
	sub_wire1(1, 102)    <= sub_wire3(102);
	sub_wire1(1, 103)    <= sub_wire3(103);
	sub_wire1(1, 104)    <= sub_wire3(104);
	sub_wire1(1, 105)    <= sub_wire3(105);
	sub_wire1(1, 106)    <= sub_wire3(106);
	sub_wire1(1, 107)    <= sub_wire3(107);
	sub_wire1(1, 108)    <= sub_wire3(108);
	sub_wire1(1, 109)    <= sub_wire3(109);
	sub_wire1(1, 110)    <= sub_wire3(110);
	sub_wire1(1, 111)    <= sub_wire3(111);
	sub_wire1(1, 112)    <= sub_wire3(112);
	sub_wire1(1, 113)    <= sub_wire3(113);
	sub_wire1(1, 114)    <= sub_wire3(114);
	sub_wire1(1, 115)    <= sub_wire3(115);
	sub_wire1(1, 116)    <= sub_wire3(116);
	sub_wire1(1, 117)    <= sub_wire3(117);
	sub_wire1(1, 118)    <= sub_wire3(118);
	sub_wire1(1, 119)    <= sub_wire3(119);
	sub_wire1(1, 120)    <= sub_wire3(120);
	sub_wire1(1, 121)    <= sub_wire3(121);
	sub_wire1(1, 122)    <= sub_wire3(122);
	sub_wire1(1, 123)    <= sub_wire3(123);
	sub_wire1(1, 124)    <= sub_wire3(124);
	sub_wire1(1, 125)    <= sub_wire3(125);
	sub_wire1(1, 126)    <= sub_wire3(126);
	sub_wire1(1, 127)    <= sub_wire3(127);
	sub_wire1(1, 128)    <= sub_wire3(128);
	sub_wire1(1, 129)    <= sub_wire3(129);
	sub_wire1(1, 130)    <= sub_wire3(130);
	sub_wire1(1, 131)    <= sub_wire3(131);
	sub_wire1(1, 132)    <= sub_wire3(132);
	sub_wire1(1, 133)    <= sub_wire3(133);
	sub_wire1(1, 134)    <= sub_wire3(134);
	sub_wire1(1, 135)    <= sub_wire3(135);
	sub_wire1(1, 136)    <= sub_wire3(136);
	sub_wire1(1, 137)    <= sub_wire3(137);
	sub_wire1(1, 138)    <= sub_wire3(138);
	sub_wire1(1, 139)    <= sub_wire3(139);
	sub_wire1(1, 140)    <= sub_wire3(140);
	sub_wire1(1, 141)    <= sub_wire3(141);
	sub_wire1(1, 142)    <= sub_wire3(142);
	sub_wire1(1, 143)    <= sub_wire3(143);
	sub_wire1(1, 144)    <= sub_wire3(144);
	sub_wire1(1, 145)    <= sub_wire3(145);
	sub_wire1(1, 146)    <= sub_wire3(146);
	sub_wire1(1, 147)    <= sub_wire3(147);
	sub_wire1(1, 148)    <= sub_wire3(148);
	sub_wire1(1, 149)    <= sub_wire3(149);
	sub_wire1(1, 150)    <= sub_wire3(150);
	sub_wire1(1, 151)    <= sub_wire3(151);
	sub_wire1(1, 152)    <= sub_wire3(152);
	sub_wire1(1, 153)    <= sub_wire3(153);
	sub_wire1(1, 154)    <= sub_wire3(154);
	sub_wire1(1, 155)    <= sub_wire3(155);
	sub_wire1(1, 156)    <= sub_wire3(156);
	sub_wire1(1, 157)    <= sub_wire3(157);
	sub_wire1(1, 158)    <= sub_wire3(158);
	sub_wire1(1, 159)    <= sub_wire3(159);
	sub_wire1(1, 160)    <= sub_wire3(160);
	sub_wire1(1, 161)    <= sub_wire3(161);
	sub_wire1(1, 162)    <= sub_wire3(162);
	sub_wire1(1, 163)    <= sub_wire3(163);
	sub_wire1(1, 164)    <= sub_wire3(164);
	sub_wire1(1, 165)    <= sub_wire3(165);
	sub_wire1(1, 166)    <= sub_wire3(166);
	sub_wire1(1, 167)    <= sub_wire3(167);
	sub_wire1(1, 168)    <= sub_wire3(168);
	sub_wire1(1, 169)    <= sub_wire3(169);
	sub_wire1(1, 170)    <= sub_wire3(170);
	sub_wire1(1, 171)    <= sub_wire3(171);
	sub_wire1(1, 172)    <= sub_wire3(172);
	sub_wire1(1, 173)    <= sub_wire3(173);
	sub_wire1(1, 174)    <= sub_wire3(174);
	sub_wire1(1, 175)    <= sub_wire3(175);
	sub_wire1(1, 176)    <= sub_wire3(176);
	sub_wire1(1, 177)    <= sub_wire3(177);
	sub_wire1(1, 178)    <= sub_wire3(178);
	sub_wire1(1, 179)    <= sub_wire3(179);
	sub_wire1(1, 180)    <= sub_wire3(180);
	sub_wire1(1, 181)    <= sub_wire3(181);
	sub_wire1(1, 182)    <= sub_wire3(182);
	sub_wire1(1, 183)    <= sub_wire3(183);
	sub_wire1(1, 184)    <= sub_wire3(184);
	sub_wire1(1, 185)    <= sub_wire3(185);
	sub_wire1(1, 186)    <= sub_wire3(186);
	sub_wire1(1, 187)    <= sub_wire3(187);
	sub_wire1(1, 188)    <= sub_wire3(188);
	sub_wire1(1, 189)    <= sub_wire3(189);
	sub_wire1(1, 190)    <= sub_wire3(190);
	sub_wire1(1, 191)    <= sub_wire3(191);
	sub_wire1(1, 192)    <= sub_wire3(192);
	sub_wire1(1, 193)    <= sub_wire3(193);
	sub_wire1(1, 194)    <= sub_wire3(194);
	sub_wire1(1, 195)    <= sub_wire3(195);
	sub_wire1(1, 196)    <= sub_wire3(196);
	sub_wire1(1, 197)    <= sub_wire3(197);
	sub_wire1(1, 198)    <= sub_wire3(198);
	sub_wire1(1, 199)    <= sub_wire3(199);
	sub_wire1(1, 200)    <= sub_wire3(200);
	sub_wire1(1, 201)    <= sub_wire3(201);
	sub_wire1(1, 202)    <= sub_wire3(202);
	sub_wire1(1, 203)    <= sub_wire3(203);
	sub_wire1(1, 204)    <= sub_wire3(204);
	sub_wire1(1, 205)    <= sub_wire3(205);
	sub_wire1(1, 206)    <= sub_wire3(206);
	sub_wire1(1, 207)    <= sub_wire3(207);
	sub_wire1(1, 208)    <= sub_wire3(208);
	sub_wire1(1, 209)    <= sub_wire3(209);
	sub_wire1(1, 210)    <= sub_wire3(210);
	sub_wire1(1, 211)    <= sub_wire3(211);
	sub_wire1(1, 212)    <= sub_wire3(212);
	sub_wire1(1, 213)    <= sub_wire3(213);
	sub_wire1(1, 214)    <= sub_wire3(214);
	sub_wire1(1, 215)    <= sub_wire3(215);
	sub_wire1(1, 216)    <= sub_wire3(216);
	sub_wire1(1, 217)    <= sub_wire3(217);
	sub_wire1(1, 218)    <= sub_wire3(218);
	sub_wire1(1, 219)    <= sub_wire3(219);
	sub_wire1(1, 220)    <= sub_wire3(220);
	sub_wire1(1, 221)    <= sub_wire3(221);
	sub_wire1(1, 222)    <= sub_wire3(222);
	sub_wire1(1, 223)    <= sub_wire3(223);
	sub_wire1(1, 224)    <= sub_wire3(224);
	sub_wire1(1, 225)    <= sub_wire3(225);
	sub_wire1(1, 226)    <= sub_wire3(226);
	sub_wire1(1, 227)    <= sub_wire3(227);
	sub_wire1(1, 228)    <= sub_wire3(228);
	sub_wire1(1, 229)    <= sub_wire3(229);
	sub_wire1(1, 230)    <= sub_wire3(230);
	sub_wire1(1, 231)    <= sub_wire3(231);
	sub_wire1(1, 232)    <= sub_wire3(232);
	sub_wire1(1, 233)    <= sub_wire3(233);
	sub_wire1(1, 234)    <= sub_wire3(234);
	sub_wire1(1, 235)    <= sub_wire3(235);
	sub_wire1(1, 236)    <= sub_wire3(236);
	sub_wire1(1, 237)    <= sub_wire3(237);
	sub_wire1(1, 238)    <= sub_wire3(238);
	sub_wire1(1, 239)    <= sub_wire3(239);
	sub_wire1(1, 240)    <= sub_wire3(240);
	sub_wire1(1, 241)    <= sub_wire3(241);
	sub_wire1(1, 242)    <= sub_wire3(242);
	sub_wire1(1, 243)    <= sub_wire3(243);
	sub_wire1(1, 244)    <= sub_wire3(244);
	sub_wire1(1, 245)    <= sub_wire3(245);
	sub_wire1(1, 246)    <= sub_wire3(246);
	sub_wire1(1, 247)    <= sub_wire3(247);
	sub_wire1(1, 248)    <= sub_wire3(248);
	sub_wire1(1, 249)    <= sub_wire3(249);
	sub_wire1(1, 250)    <= sub_wire3(250);
	sub_wire1(1, 251)    <= sub_wire3(251);
	sub_wire1(1, 252)    <= sub_wire3(252);
	sub_wire1(1, 253)    <= sub_wire3(253);
	sub_wire1(1, 254)    <= sub_wire3(254);
	sub_wire1(1, 255)    <= sub_wire3(255);
	sub_wire1(0, 0)    <= sub_wire4(0);
	sub_wire1(0, 1)    <= sub_wire4(1);
	sub_wire1(0, 2)    <= sub_wire4(2);
	sub_wire1(0, 3)    <= sub_wire4(3);
	sub_wire1(0, 4)    <= sub_wire4(4);
	sub_wire1(0, 5)    <= sub_wire4(5);
	sub_wire1(0, 6)    <= sub_wire4(6);
	sub_wire1(0, 7)    <= sub_wire4(7);
	sub_wire1(0, 8)    <= sub_wire4(8);
	sub_wire1(0, 9)    <= sub_wire4(9);
	sub_wire1(0, 10)    <= sub_wire4(10);
	sub_wire1(0, 11)    <= sub_wire4(11);
	sub_wire1(0, 12)    <= sub_wire4(12);
	sub_wire1(0, 13)    <= sub_wire4(13);
	sub_wire1(0, 14)    <= sub_wire4(14);
	sub_wire1(0, 15)    <= sub_wire4(15);
	sub_wire1(0, 16)    <= sub_wire4(16);
	sub_wire1(0, 17)    <= sub_wire4(17);
	sub_wire1(0, 18)    <= sub_wire4(18);
	sub_wire1(0, 19)    <= sub_wire4(19);
	sub_wire1(0, 20)    <= sub_wire4(20);
	sub_wire1(0, 21)    <= sub_wire4(21);
	sub_wire1(0, 22)    <= sub_wire4(22);
	sub_wire1(0, 23)    <= sub_wire4(23);
	sub_wire1(0, 24)    <= sub_wire4(24);
	sub_wire1(0, 25)    <= sub_wire4(25);
	sub_wire1(0, 26)    <= sub_wire4(26);
	sub_wire1(0, 27)    <= sub_wire4(27);
	sub_wire1(0, 28)    <= sub_wire4(28);
	sub_wire1(0, 29)    <= sub_wire4(29);
	sub_wire1(0, 30)    <= sub_wire4(30);
	sub_wire1(0, 31)    <= sub_wire4(31);
	sub_wire1(0, 32)    <= sub_wire4(32);
	sub_wire1(0, 33)    <= sub_wire4(33);
	sub_wire1(0, 34)    <= sub_wire4(34);
	sub_wire1(0, 35)    <= sub_wire4(35);
	sub_wire1(0, 36)    <= sub_wire4(36);
	sub_wire1(0, 37)    <= sub_wire4(37);
	sub_wire1(0, 38)    <= sub_wire4(38);
	sub_wire1(0, 39)    <= sub_wire4(39);
	sub_wire1(0, 40)    <= sub_wire4(40);
	sub_wire1(0, 41)    <= sub_wire4(41);
	sub_wire1(0, 42)    <= sub_wire4(42);
	sub_wire1(0, 43)    <= sub_wire4(43);
	sub_wire1(0, 44)    <= sub_wire4(44);
	sub_wire1(0, 45)    <= sub_wire4(45);
	sub_wire1(0, 46)    <= sub_wire4(46);
	sub_wire1(0, 47)    <= sub_wire4(47);
	sub_wire1(0, 48)    <= sub_wire4(48);
	sub_wire1(0, 49)    <= sub_wire4(49);
	sub_wire1(0, 50)    <= sub_wire4(50);
	sub_wire1(0, 51)    <= sub_wire4(51);
	sub_wire1(0, 52)    <= sub_wire4(52);
	sub_wire1(0, 53)    <= sub_wire4(53);
	sub_wire1(0, 54)    <= sub_wire4(54);
	sub_wire1(0, 55)    <= sub_wire4(55);
	sub_wire1(0, 56)    <= sub_wire4(56);
	sub_wire1(0, 57)    <= sub_wire4(57);
	sub_wire1(0, 58)    <= sub_wire4(58);
	sub_wire1(0, 59)    <= sub_wire4(59);
	sub_wire1(0, 60)    <= sub_wire4(60);
	sub_wire1(0, 61)    <= sub_wire4(61);
	sub_wire1(0, 62)    <= sub_wire4(62);
	sub_wire1(0, 63)    <= sub_wire4(63);
	sub_wire1(0, 64)    <= sub_wire4(64);
	sub_wire1(0, 65)    <= sub_wire4(65);
	sub_wire1(0, 66)    <= sub_wire4(66);
	sub_wire1(0, 67)    <= sub_wire4(67);
	sub_wire1(0, 68)    <= sub_wire4(68);
	sub_wire1(0, 69)    <= sub_wire4(69);
	sub_wire1(0, 70)    <= sub_wire4(70);
	sub_wire1(0, 71)    <= sub_wire4(71);
	sub_wire1(0, 72)    <= sub_wire4(72);
	sub_wire1(0, 73)    <= sub_wire4(73);
	sub_wire1(0, 74)    <= sub_wire4(74);
	sub_wire1(0, 75)    <= sub_wire4(75);
	sub_wire1(0, 76)    <= sub_wire4(76);
	sub_wire1(0, 77)    <= sub_wire4(77);
	sub_wire1(0, 78)    <= sub_wire4(78);
	sub_wire1(0, 79)    <= sub_wire4(79);
	sub_wire1(0, 80)    <= sub_wire4(80);
	sub_wire1(0, 81)    <= sub_wire4(81);
	sub_wire1(0, 82)    <= sub_wire4(82);
	sub_wire1(0, 83)    <= sub_wire4(83);
	sub_wire1(0, 84)    <= sub_wire4(84);
	sub_wire1(0, 85)    <= sub_wire4(85);
	sub_wire1(0, 86)    <= sub_wire4(86);
	sub_wire1(0, 87)    <= sub_wire4(87);
	sub_wire1(0, 88)    <= sub_wire4(88);
	sub_wire1(0, 89)    <= sub_wire4(89);
	sub_wire1(0, 90)    <= sub_wire4(90);
	sub_wire1(0, 91)    <= sub_wire4(91);
	sub_wire1(0, 92)    <= sub_wire4(92);
	sub_wire1(0, 93)    <= sub_wire4(93);
	sub_wire1(0, 94)    <= sub_wire4(94);
	sub_wire1(0, 95)    <= sub_wire4(95);
	sub_wire1(0, 96)    <= sub_wire4(96);
	sub_wire1(0, 97)    <= sub_wire4(97);
	sub_wire1(0, 98)    <= sub_wire4(98);
	sub_wire1(0, 99)    <= sub_wire4(99);
	sub_wire1(0, 100)    <= sub_wire4(100);
	sub_wire1(0, 101)    <= sub_wire4(101);
	sub_wire1(0, 102)    <= sub_wire4(102);
	sub_wire1(0, 103)    <= sub_wire4(103);
	sub_wire1(0, 104)    <= sub_wire4(104);
	sub_wire1(0, 105)    <= sub_wire4(105);
	sub_wire1(0, 106)    <= sub_wire4(106);
	sub_wire1(0, 107)    <= sub_wire4(107);
	sub_wire1(0, 108)    <= sub_wire4(108);
	sub_wire1(0, 109)    <= sub_wire4(109);
	sub_wire1(0, 110)    <= sub_wire4(110);
	sub_wire1(0, 111)    <= sub_wire4(111);
	sub_wire1(0, 112)    <= sub_wire4(112);
	sub_wire1(0, 113)    <= sub_wire4(113);
	sub_wire1(0, 114)    <= sub_wire4(114);
	sub_wire1(0, 115)    <= sub_wire4(115);
	sub_wire1(0, 116)    <= sub_wire4(116);
	sub_wire1(0, 117)    <= sub_wire4(117);
	sub_wire1(0, 118)    <= sub_wire4(118);
	sub_wire1(0, 119)    <= sub_wire4(119);
	sub_wire1(0, 120)    <= sub_wire4(120);
	sub_wire1(0, 121)    <= sub_wire4(121);
	sub_wire1(0, 122)    <= sub_wire4(122);
	sub_wire1(0, 123)    <= sub_wire4(123);
	sub_wire1(0, 124)    <= sub_wire4(124);
	sub_wire1(0, 125)    <= sub_wire4(125);
	sub_wire1(0, 126)    <= sub_wire4(126);
	sub_wire1(0, 127)    <= sub_wire4(127);
	sub_wire1(0, 128)    <= sub_wire4(128);
	sub_wire1(0, 129)    <= sub_wire4(129);
	sub_wire1(0, 130)    <= sub_wire4(130);
	sub_wire1(0, 131)    <= sub_wire4(131);
	sub_wire1(0, 132)    <= sub_wire4(132);
	sub_wire1(0, 133)    <= sub_wire4(133);
	sub_wire1(0, 134)    <= sub_wire4(134);
	sub_wire1(0, 135)    <= sub_wire4(135);
	sub_wire1(0, 136)    <= sub_wire4(136);
	sub_wire1(0, 137)    <= sub_wire4(137);
	sub_wire1(0, 138)    <= sub_wire4(138);
	sub_wire1(0, 139)    <= sub_wire4(139);
	sub_wire1(0, 140)    <= sub_wire4(140);
	sub_wire1(0, 141)    <= sub_wire4(141);
	sub_wire1(0, 142)    <= sub_wire4(142);
	sub_wire1(0, 143)    <= sub_wire4(143);
	sub_wire1(0, 144)    <= sub_wire4(144);
	sub_wire1(0, 145)    <= sub_wire4(145);
	sub_wire1(0, 146)    <= sub_wire4(146);
	sub_wire1(0, 147)    <= sub_wire4(147);
	sub_wire1(0, 148)    <= sub_wire4(148);
	sub_wire1(0, 149)    <= sub_wire4(149);
	sub_wire1(0, 150)    <= sub_wire4(150);
	sub_wire1(0, 151)    <= sub_wire4(151);
	sub_wire1(0, 152)    <= sub_wire4(152);
	sub_wire1(0, 153)    <= sub_wire4(153);
	sub_wire1(0, 154)    <= sub_wire4(154);
	sub_wire1(0, 155)    <= sub_wire4(155);
	sub_wire1(0, 156)    <= sub_wire4(156);
	sub_wire1(0, 157)    <= sub_wire4(157);
	sub_wire1(0, 158)    <= sub_wire4(158);
	sub_wire1(0, 159)    <= sub_wire4(159);
	sub_wire1(0, 160)    <= sub_wire4(160);
	sub_wire1(0, 161)    <= sub_wire4(161);
	sub_wire1(0, 162)    <= sub_wire4(162);
	sub_wire1(0, 163)    <= sub_wire4(163);
	sub_wire1(0, 164)    <= sub_wire4(164);
	sub_wire1(0, 165)    <= sub_wire4(165);
	sub_wire1(0, 166)    <= sub_wire4(166);
	sub_wire1(0, 167)    <= sub_wire4(167);
	sub_wire1(0, 168)    <= sub_wire4(168);
	sub_wire1(0, 169)    <= sub_wire4(169);
	sub_wire1(0, 170)    <= sub_wire4(170);
	sub_wire1(0, 171)    <= sub_wire4(171);
	sub_wire1(0, 172)    <= sub_wire4(172);
	sub_wire1(0, 173)    <= sub_wire4(173);
	sub_wire1(0, 174)    <= sub_wire4(174);
	sub_wire1(0, 175)    <= sub_wire4(175);
	sub_wire1(0, 176)    <= sub_wire4(176);
	sub_wire1(0, 177)    <= sub_wire4(177);
	sub_wire1(0, 178)    <= sub_wire4(178);
	sub_wire1(0, 179)    <= sub_wire4(179);
	sub_wire1(0, 180)    <= sub_wire4(180);
	sub_wire1(0, 181)    <= sub_wire4(181);
	sub_wire1(0, 182)    <= sub_wire4(182);
	sub_wire1(0, 183)    <= sub_wire4(183);
	sub_wire1(0, 184)    <= sub_wire4(184);
	sub_wire1(0, 185)    <= sub_wire4(185);
	sub_wire1(0, 186)    <= sub_wire4(186);
	sub_wire1(0, 187)    <= sub_wire4(187);
	sub_wire1(0, 188)    <= sub_wire4(188);
	sub_wire1(0, 189)    <= sub_wire4(189);
	sub_wire1(0, 190)    <= sub_wire4(190);
	sub_wire1(0, 191)    <= sub_wire4(191);
	sub_wire1(0, 192)    <= sub_wire4(192);
	sub_wire1(0, 193)    <= sub_wire4(193);
	sub_wire1(0, 194)    <= sub_wire4(194);
	sub_wire1(0, 195)    <= sub_wire4(195);
	sub_wire1(0, 196)    <= sub_wire4(196);
	sub_wire1(0, 197)    <= sub_wire4(197);
	sub_wire1(0, 198)    <= sub_wire4(198);
	sub_wire1(0, 199)    <= sub_wire4(199);
	sub_wire1(0, 200)    <= sub_wire4(200);
	sub_wire1(0, 201)    <= sub_wire4(201);
	sub_wire1(0, 202)    <= sub_wire4(202);
	sub_wire1(0, 203)    <= sub_wire4(203);
	sub_wire1(0, 204)    <= sub_wire4(204);
	sub_wire1(0, 205)    <= sub_wire4(205);
	sub_wire1(0, 206)    <= sub_wire4(206);
	sub_wire1(0, 207)    <= sub_wire4(207);
	sub_wire1(0, 208)    <= sub_wire4(208);
	sub_wire1(0, 209)    <= sub_wire4(209);
	sub_wire1(0, 210)    <= sub_wire4(210);
	sub_wire1(0, 211)    <= sub_wire4(211);
	sub_wire1(0, 212)    <= sub_wire4(212);
	sub_wire1(0, 213)    <= sub_wire4(213);
	sub_wire1(0, 214)    <= sub_wire4(214);
	sub_wire1(0, 215)    <= sub_wire4(215);
	sub_wire1(0, 216)    <= sub_wire4(216);
	sub_wire1(0, 217)    <= sub_wire4(217);
	sub_wire1(0, 218)    <= sub_wire4(218);
	sub_wire1(0, 219)    <= sub_wire4(219);
	sub_wire1(0, 220)    <= sub_wire4(220);
	sub_wire1(0, 221)    <= sub_wire4(221);
	sub_wire1(0, 222)    <= sub_wire4(222);
	sub_wire1(0, 223)    <= sub_wire4(223);
	sub_wire1(0, 224)    <= sub_wire4(224);
	sub_wire1(0, 225)    <= sub_wire4(225);
	sub_wire1(0, 226)    <= sub_wire4(226);
	sub_wire1(0, 227)    <= sub_wire4(227);
	sub_wire1(0, 228)    <= sub_wire4(228);
	sub_wire1(0, 229)    <= sub_wire4(229);
	sub_wire1(0, 230)    <= sub_wire4(230);
	sub_wire1(0, 231)    <= sub_wire4(231);
	sub_wire1(0, 232)    <= sub_wire4(232);
	sub_wire1(0, 233)    <= sub_wire4(233);
	sub_wire1(0, 234)    <= sub_wire4(234);
	sub_wire1(0, 235)    <= sub_wire4(235);
	sub_wire1(0, 236)    <= sub_wire4(236);
	sub_wire1(0, 237)    <= sub_wire4(237);
	sub_wire1(0, 238)    <= sub_wire4(238);
	sub_wire1(0, 239)    <= sub_wire4(239);
	sub_wire1(0, 240)    <= sub_wire4(240);
	sub_wire1(0, 241)    <= sub_wire4(241);
	sub_wire1(0, 242)    <= sub_wire4(242);
	sub_wire1(0, 243)    <= sub_wire4(243);
	sub_wire1(0, 244)    <= sub_wire4(244);
	sub_wire1(0, 245)    <= sub_wire4(245);
	sub_wire1(0, 246)    <= sub_wire4(246);
	sub_wire1(0, 247)    <= sub_wire4(247);
	sub_wire1(0, 248)    <= sub_wire4(248);
	sub_wire1(0, 249)    <= sub_wire4(249);
	sub_wire1(0, 250)    <= sub_wire4(250);
	sub_wire1(0, 251)    <= sub_wire4(251);
	sub_wire1(0, 252)    <= sub_wire4(252);
	sub_wire1(0, 253)    <= sub_wire4(253);
	sub_wire1(0, 254)    <= sub_wire4(254);
	sub_wire1(0, 255)    <= sub_wire4(255);
	result    <= sub_wire5(255 DOWNTO 0);

	LPM_MUX_component : LPM_MUX
	GENERIC MAP (
		lpm_pipeline => 1,
		lpm_size => 4,
		lpm_type => "LPM_MUX",
		lpm_width => 256,
		lpm_widths => 2
	)
	PORT MAP (
		clock => clock,
		data => sub_wire1,
		sel => sel,
		result => sub_wire5
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "1"
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "4"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "256"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "2"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data0x 0 0 256 0 INPUT NODEFVAL "data0x[255..0]"
-- Retrieval info: USED_PORT: data1x 0 0 256 0 INPUT NODEFVAL "data1x[255..0]"
-- Retrieval info: USED_PORT: data2x 0 0 256 0 INPUT NODEFVAL "data2x[255..0]"
-- Retrieval info: USED_PORT: data3x 0 0 256 0 INPUT NODEFVAL "data3x[255..0]"
-- Retrieval info: USED_PORT: result 0 0 256 0 OUTPUT NODEFVAL "result[255..0]"
-- Retrieval info: USED_PORT: sel 0 0 2 0 INPUT NODEFVAL "sel[1..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data 1 0 256 0 data0x 0 0 256 0
-- Retrieval info: CONNECT: @data 1 1 256 0 data1x 0 0 256 0
-- Retrieval info: CONNECT: @data 1 2 256 0 data2x 0 0 256 0
-- Retrieval info: CONNECT: @data 1 3 256 0 data3x 0 0 256 0
-- Retrieval info: CONNECT: @sel 0 0 2 0 sel 0 0 2 0
-- Retrieval info: CONNECT: result 0 0 256 0 @result 0 0 256 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX4_256b.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX4_256b.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX4_256b.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX4_256b.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX4_256b_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
