-- megafunction wizard: %PARALLEL_ADD%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: parallel_add 

-- ============================================================
-- File Name: Turn_Adder.vhd
-- Megafunction Name(s):
-- 			parallel_add
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 15.0.0 Build 145 04/22/2015 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus II License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY Turn_Adder IS
	PORT
	(
		aclr		: IN STD_LOGIC  := '0';
		clock		: IN STD_LOGIC  := '0';
		data0x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data10x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data11x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data12x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data13x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data14x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data15x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data16x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data17x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data18x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data19x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data20x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data21x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data22x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data23x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data24x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data25x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data26x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data27x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data28x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data29x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data30x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data31x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data32x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data33x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data34x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data35x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data36x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data8x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		data9x		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (14 DOWNTO 0)
	);
END Turn_Adder;


ARCHITECTURE SYN OF turn_adder IS

--	type ALTERA_MF_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire1	: ALTERA_MF_LOGIC_2D (36 DOWNTO 0, 8 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire14	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire15	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire16	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire17	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire18	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire19	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire20	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire21	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire22	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire23	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire24	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire25	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire26	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire27	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire28	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire29	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire30	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire31	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire32	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire33	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire34	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire35	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire36	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire37	: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL sub_wire38	: STD_LOGIC_VECTOR (14 DOWNTO 0);

BEGIN
	sub_wire37    <= data0x(8 DOWNTO 0);
	sub_wire36    <= data1x(8 DOWNTO 0);
	sub_wire35    <= data2x(8 DOWNTO 0);
	sub_wire34    <= data3x(8 DOWNTO 0);
	sub_wire33    <= data4x(8 DOWNTO 0);
	sub_wire32    <= data5x(8 DOWNTO 0);
	sub_wire31    <= data6x(8 DOWNTO 0);
	sub_wire30    <= data7x(8 DOWNTO 0);
	sub_wire29    <= data8x(8 DOWNTO 0);
	sub_wire28    <= data9x(8 DOWNTO 0);
	sub_wire27    <= data10x(8 DOWNTO 0);
	sub_wire26    <= data11x(8 DOWNTO 0);
	sub_wire25    <= data12x(8 DOWNTO 0);
	sub_wire24    <= data13x(8 DOWNTO 0);
	sub_wire23    <= data14x(8 DOWNTO 0);
	sub_wire22    <= data15x(8 DOWNTO 0);
	sub_wire21    <= data16x(8 DOWNTO 0);
	sub_wire20    <= data17x(8 DOWNTO 0);
	sub_wire19    <= data18x(8 DOWNTO 0);
	sub_wire18    <= data19x(8 DOWNTO 0);
	sub_wire17    <= data20x(8 DOWNTO 0);
	sub_wire16    <= data21x(8 DOWNTO 0);
	sub_wire15    <= data22x(8 DOWNTO 0);
	sub_wire14    <= data23x(8 DOWNTO 0);
	sub_wire13    <= data24x(8 DOWNTO 0);
	sub_wire12    <= data25x(8 DOWNTO 0);
	sub_wire11    <= data26x(8 DOWNTO 0);
	sub_wire10    <= data27x(8 DOWNTO 0);
	sub_wire9    <= data28x(8 DOWNTO 0);
	sub_wire8    <= data29x(8 DOWNTO 0);
	sub_wire7    <= data30x(8 DOWNTO 0);
	sub_wire6    <= data31x(8 DOWNTO 0);
	sub_wire5    <= data32x(8 DOWNTO 0);
	sub_wire4    <= data33x(8 DOWNTO 0);
	sub_wire3    <= data34x(8 DOWNTO 0);
	sub_wire2    <= data35x(8 DOWNTO 0);
	sub_wire0    <= data36x(8 DOWNTO 0);
	sub_wire1(36, 0)    <= sub_wire0(0);
	sub_wire1(36, 1)    <= sub_wire0(1);
	sub_wire1(36, 2)    <= sub_wire0(2);
	sub_wire1(36, 3)    <= sub_wire0(3);
	sub_wire1(36, 4)    <= sub_wire0(4);
	sub_wire1(36, 5)    <= sub_wire0(5);
	sub_wire1(36, 6)    <= sub_wire0(6);
	sub_wire1(36, 7)    <= sub_wire0(7);
	sub_wire1(36, 8)    <= sub_wire0(8);
	sub_wire1(35, 0)    <= sub_wire2(0);
	sub_wire1(35, 1)    <= sub_wire2(1);
	sub_wire1(35, 2)    <= sub_wire2(2);
	sub_wire1(35, 3)    <= sub_wire2(3);
	sub_wire1(35, 4)    <= sub_wire2(4);
	sub_wire1(35, 5)    <= sub_wire2(5);
	sub_wire1(35, 6)    <= sub_wire2(6);
	sub_wire1(35, 7)    <= sub_wire2(7);
	sub_wire1(35, 8)    <= sub_wire2(8);
	sub_wire1(34, 0)    <= sub_wire3(0);
	sub_wire1(34, 1)    <= sub_wire3(1);
	sub_wire1(34, 2)    <= sub_wire3(2);
	sub_wire1(34, 3)    <= sub_wire3(3);
	sub_wire1(34, 4)    <= sub_wire3(4);
	sub_wire1(34, 5)    <= sub_wire3(5);
	sub_wire1(34, 6)    <= sub_wire3(6);
	sub_wire1(34, 7)    <= sub_wire3(7);
	sub_wire1(34, 8)    <= sub_wire3(8);
	sub_wire1(33, 0)    <= sub_wire4(0);
	sub_wire1(33, 1)    <= sub_wire4(1);
	sub_wire1(33, 2)    <= sub_wire4(2);
	sub_wire1(33, 3)    <= sub_wire4(3);
	sub_wire1(33, 4)    <= sub_wire4(4);
	sub_wire1(33, 5)    <= sub_wire4(5);
	sub_wire1(33, 6)    <= sub_wire4(6);
	sub_wire1(33, 7)    <= sub_wire4(7);
	sub_wire1(33, 8)    <= sub_wire4(8);
	sub_wire1(32, 0)    <= sub_wire5(0);
	sub_wire1(32, 1)    <= sub_wire5(1);
	sub_wire1(32, 2)    <= sub_wire5(2);
	sub_wire1(32, 3)    <= sub_wire5(3);
	sub_wire1(32, 4)    <= sub_wire5(4);
	sub_wire1(32, 5)    <= sub_wire5(5);
	sub_wire1(32, 6)    <= sub_wire5(6);
	sub_wire1(32, 7)    <= sub_wire5(7);
	sub_wire1(32, 8)    <= sub_wire5(8);
	sub_wire1(31, 0)    <= sub_wire6(0);
	sub_wire1(31, 1)    <= sub_wire6(1);
	sub_wire1(31, 2)    <= sub_wire6(2);
	sub_wire1(31, 3)    <= sub_wire6(3);
	sub_wire1(31, 4)    <= sub_wire6(4);
	sub_wire1(31, 5)    <= sub_wire6(5);
	sub_wire1(31, 6)    <= sub_wire6(6);
	sub_wire1(31, 7)    <= sub_wire6(7);
	sub_wire1(31, 8)    <= sub_wire6(8);
	sub_wire1(30, 0)    <= sub_wire7(0);
	sub_wire1(30, 1)    <= sub_wire7(1);
	sub_wire1(30, 2)    <= sub_wire7(2);
	sub_wire1(30, 3)    <= sub_wire7(3);
	sub_wire1(30, 4)    <= sub_wire7(4);
	sub_wire1(30, 5)    <= sub_wire7(5);
	sub_wire1(30, 6)    <= sub_wire7(6);
	sub_wire1(30, 7)    <= sub_wire7(7);
	sub_wire1(30, 8)    <= sub_wire7(8);
	sub_wire1(29, 0)    <= sub_wire8(0);
	sub_wire1(29, 1)    <= sub_wire8(1);
	sub_wire1(29, 2)    <= sub_wire8(2);
	sub_wire1(29, 3)    <= sub_wire8(3);
	sub_wire1(29, 4)    <= sub_wire8(4);
	sub_wire1(29, 5)    <= sub_wire8(5);
	sub_wire1(29, 6)    <= sub_wire8(6);
	sub_wire1(29, 7)    <= sub_wire8(7);
	sub_wire1(29, 8)    <= sub_wire8(8);
	sub_wire1(28, 0)    <= sub_wire9(0);
	sub_wire1(28, 1)    <= sub_wire9(1);
	sub_wire1(28, 2)    <= sub_wire9(2);
	sub_wire1(28, 3)    <= sub_wire9(3);
	sub_wire1(28, 4)    <= sub_wire9(4);
	sub_wire1(28, 5)    <= sub_wire9(5);
	sub_wire1(28, 6)    <= sub_wire9(6);
	sub_wire1(28, 7)    <= sub_wire9(7);
	sub_wire1(28, 8)    <= sub_wire9(8);
	sub_wire1(27, 0)    <= sub_wire10(0);
	sub_wire1(27, 1)    <= sub_wire10(1);
	sub_wire1(27, 2)    <= sub_wire10(2);
	sub_wire1(27, 3)    <= sub_wire10(3);
	sub_wire1(27, 4)    <= sub_wire10(4);
	sub_wire1(27, 5)    <= sub_wire10(5);
	sub_wire1(27, 6)    <= sub_wire10(6);
	sub_wire1(27, 7)    <= sub_wire10(7);
	sub_wire1(27, 8)    <= sub_wire10(8);
	sub_wire1(26, 0)    <= sub_wire11(0);
	sub_wire1(26, 1)    <= sub_wire11(1);
	sub_wire1(26, 2)    <= sub_wire11(2);
	sub_wire1(26, 3)    <= sub_wire11(3);
	sub_wire1(26, 4)    <= sub_wire11(4);
	sub_wire1(26, 5)    <= sub_wire11(5);
	sub_wire1(26, 6)    <= sub_wire11(6);
	sub_wire1(26, 7)    <= sub_wire11(7);
	sub_wire1(26, 8)    <= sub_wire11(8);
	sub_wire1(25, 0)    <= sub_wire12(0);
	sub_wire1(25, 1)    <= sub_wire12(1);
	sub_wire1(25, 2)    <= sub_wire12(2);
	sub_wire1(25, 3)    <= sub_wire12(3);
	sub_wire1(25, 4)    <= sub_wire12(4);
	sub_wire1(25, 5)    <= sub_wire12(5);
	sub_wire1(25, 6)    <= sub_wire12(6);
	sub_wire1(25, 7)    <= sub_wire12(7);
	sub_wire1(25, 8)    <= sub_wire12(8);
	sub_wire1(24, 0)    <= sub_wire13(0);
	sub_wire1(24, 1)    <= sub_wire13(1);
	sub_wire1(24, 2)    <= sub_wire13(2);
	sub_wire1(24, 3)    <= sub_wire13(3);
	sub_wire1(24, 4)    <= sub_wire13(4);
	sub_wire1(24, 5)    <= sub_wire13(5);
	sub_wire1(24, 6)    <= sub_wire13(6);
	sub_wire1(24, 7)    <= sub_wire13(7);
	sub_wire1(24, 8)    <= sub_wire13(8);
	sub_wire1(23, 0)    <= sub_wire14(0);
	sub_wire1(23, 1)    <= sub_wire14(1);
	sub_wire1(23, 2)    <= sub_wire14(2);
	sub_wire1(23, 3)    <= sub_wire14(3);
	sub_wire1(23, 4)    <= sub_wire14(4);
	sub_wire1(23, 5)    <= sub_wire14(5);
	sub_wire1(23, 6)    <= sub_wire14(6);
	sub_wire1(23, 7)    <= sub_wire14(7);
	sub_wire1(23, 8)    <= sub_wire14(8);
	sub_wire1(22, 0)    <= sub_wire15(0);
	sub_wire1(22, 1)    <= sub_wire15(1);
	sub_wire1(22, 2)    <= sub_wire15(2);
	sub_wire1(22, 3)    <= sub_wire15(3);
	sub_wire1(22, 4)    <= sub_wire15(4);
	sub_wire1(22, 5)    <= sub_wire15(5);
	sub_wire1(22, 6)    <= sub_wire15(6);
	sub_wire1(22, 7)    <= sub_wire15(7);
	sub_wire1(22, 8)    <= sub_wire15(8);
	sub_wire1(21, 0)    <= sub_wire16(0);
	sub_wire1(21, 1)    <= sub_wire16(1);
	sub_wire1(21, 2)    <= sub_wire16(2);
	sub_wire1(21, 3)    <= sub_wire16(3);
	sub_wire1(21, 4)    <= sub_wire16(4);
	sub_wire1(21, 5)    <= sub_wire16(5);
	sub_wire1(21, 6)    <= sub_wire16(6);
	sub_wire1(21, 7)    <= sub_wire16(7);
	sub_wire1(21, 8)    <= sub_wire16(8);
	sub_wire1(20, 0)    <= sub_wire17(0);
	sub_wire1(20, 1)    <= sub_wire17(1);
	sub_wire1(20, 2)    <= sub_wire17(2);
	sub_wire1(20, 3)    <= sub_wire17(3);
	sub_wire1(20, 4)    <= sub_wire17(4);
	sub_wire1(20, 5)    <= sub_wire17(5);
	sub_wire1(20, 6)    <= sub_wire17(6);
	sub_wire1(20, 7)    <= sub_wire17(7);
	sub_wire1(20, 8)    <= sub_wire17(8);
	sub_wire1(19, 0)    <= sub_wire18(0);
	sub_wire1(19, 1)    <= sub_wire18(1);
	sub_wire1(19, 2)    <= sub_wire18(2);
	sub_wire1(19, 3)    <= sub_wire18(3);
	sub_wire1(19, 4)    <= sub_wire18(4);
	sub_wire1(19, 5)    <= sub_wire18(5);
	sub_wire1(19, 6)    <= sub_wire18(6);
	sub_wire1(19, 7)    <= sub_wire18(7);
	sub_wire1(19, 8)    <= sub_wire18(8);
	sub_wire1(18, 0)    <= sub_wire19(0);
	sub_wire1(18, 1)    <= sub_wire19(1);
	sub_wire1(18, 2)    <= sub_wire19(2);
	sub_wire1(18, 3)    <= sub_wire19(3);
	sub_wire1(18, 4)    <= sub_wire19(4);
	sub_wire1(18, 5)    <= sub_wire19(5);
	sub_wire1(18, 6)    <= sub_wire19(6);
	sub_wire1(18, 7)    <= sub_wire19(7);
	sub_wire1(18, 8)    <= sub_wire19(8);
	sub_wire1(17, 0)    <= sub_wire20(0);
	sub_wire1(17, 1)    <= sub_wire20(1);
	sub_wire1(17, 2)    <= sub_wire20(2);
	sub_wire1(17, 3)    <= sub_wire20(3);
	sub_wire1(17, 4)    <= sub_wire20(4);
	sub_wire1(17, 5)    <= sub_wire20(5);
	sub_wire1(17, 6)    <= sub_wire20(6);
	sub_wire1(17, 7)    <= sub_wire20(7);
	sub_wire1(17, 8)    <= sub_wire20(8);
	sub_wire1(16, 0)    <= sub_wire21(0);
	sub_wire1(16, 1)    <= sub_wire21(1);
	sub_wire1(16, 2)    <= sub_wire21(2);
	sub_wire1(16, 3)    <= sub_wire21(3);
	sub_wire1(16, 4)    <= sub_wire21(4);
	sub_wire1(16, 5)    <= sub_wire21(5);
	sub_wire1(16, 6)    <= sub_wire21(6);
	sub_wire1(16, 7)    <= sub_wire21(7);
	sub_wire1(16, 8)    <= sub_wire21(8);
	sub_wire1(15, 0)    <= sub_wire22(0);
	sub_wire1(15, 1)    <= sub_wire22(1);
	sub_wire1(15, 2)    <= sub_wire22(2);
	sub_wire1(15, 3)    <= sub_wire22(3);
	sub_wire1(15, 4)    <= sub_wire22(4);
	sub_wire1(15, 5)    <= sub_wire22(5);
	sub_wire1(15, 6)    <= sub_wire22(6);
	sub_wire1(15, 7)    <= sub_wire22(7);
	sub_wire1(15, 8)    <= sub_wire22(8);
	sub_wire1(14, 0)    <= sub_wire23(0);
	sub_wire1(14, 1)    <= sub_wire23(1);
	sub_wire1(14, 2)    <= sub_wire23(2);
	sub_wire1(14, 3)    <= sub_wire23(3);
	sub_wire1(14, 4)    <= sub_wire23(4);
	sub_wire1(14, 5)    <= sub_wire23(5);
	sub_wire1(14, 6)    <= sub_wire23(6);
	sub_wire1(14, 7)    <= sub_wire23(7);
	sub_wire1(14, 8)    <= sub_wire23(8);
	sub_wire1(13, 0)    <= sub_wire24(0);
	sub_wire1(13, 1)    <= sub_wire24(1);
	sub_wire1(13, 2)    <= sub_wire24(2);
	sub_wire1(13, 3)    <= sub_wire24(3);
	sub_wire1(13, 4)    <= sub_wire24(4);
	sub_wire1(13, 5)    <= sub_wire24(5);
	sub_wire1(13, 6)    <= sub_wire24(6);
	sub_wire1(13, 7)    <= sub_wire24(7);
	sub_wire1(13, 8)    <= sub_wire24(8);
	sub_wire1(12, 0)    <= sub_wire25(0);
	sub_wire1(12, 1)    <= sub_wire25(1);
	sub_wire1(12, 2)    <= sub_wire25(2);
	sub_wire1(12, 3)    <= sub_wire25(3);
	sub_wire1(12, 4)    <= sub_wire25(4);
	sub_wire1(12, 5)    <= sub_wire25(5);
	sub_wire1(12, 6)    <= sub_wire25(6);
	sub_wire1(12, 7)    <= sub_wire25(7);
	sub_wire1(12, 8)    <= sub_wire25(8);
	sub_wire1(11, 0)    <= sub_wire26(0);
	sub_wire1(11, 1)    <= sub_wire26(1);
	sub_wire1(11, 2)    <= sub_wire26(2);
	sub_wire1(11, 3)    <= sub_wire26(3);
	sub_wire1(11, 4)    <= sub_wire26(4);
	sub_wire1(11, 5)    <= sub_wire26(5);
	sub_wire1(11, 6)    <= sub_wire26(6);
	sub_wire1(11, 7)    <= sub_wire26(7);
	sub_wire1(11, 8)    <= sub_wire26(8);
	sub_wire1(10, 0)    <= sub_wire27(0);
	sub_wire1(10, 1)    <= sub_wire27(1);
	sub_wire1(10, 2)    <= sub_wire27(2);
	sub_wire1(10, 3)    <= sub_wire27(3);
	sub_wire1(10, 4)    <= sub_wire27(4);
	sub_wire1(10, 5)    <= sub_wire27(5);
	sub_wire1(10, 6)    <= sub_wire27(6);
	sub_wire1(10, 7)    <= sub_wire27(7);
	sub_wire1(10, 8)    <= sub_wire27(8);
	sub_wire1(9, 0)    <= sub_wire28(0);
	sub_wire1(9, 1)    <= sub_wire28(1);
	sub_wire1(9, 2)    <= sub_wire28(2);
	sub_wire1(9, 3)    <= sub_wire28(3);
	sub_wire1(9, 4)    <= sub_wire28(4);
	sub_wire1(9, 5)    <= sub_wire28(5);
	sub_wire1(9, 6)    <= sub_wire28(6);
	sub_wire1(9, 7)    <= sub_wire28(7);
	sub_wire1(9, 8)    <= sub_wire28(8);
	sub_wire1(8, 0)    <= sub_wire29(0);
	sub_wire1(8, 1)    <= sub_wire29(1);
	sub_wire1(8, 2)    <= sub_wire29(2);
	sub_wire1(8, 3)    <= sub_wire29(3);
	sub_wire1(8, 4)    <= sub_wire29(4);
	sub_wire1(8, 5)    <= sub_wire29(5);
	sub_wire1(8, 6)    <= sub_wire29(6);
	sub_wire1(8, 7)    <= sub_wire29(7);
	sub_wire1(8, 8)    <= sub_wire29(8);
	sub_wire1(7, 0)    <= sub_wire30(0);
	sub_wire1(7, 1)    <= sub_wire30(1);
	sub_wire1(7, 2)    <= sub_wire30(2);
	sub_wire1(7, 3)    <= sub_wire30(3);
	sub_wire1(7, 4)    <= sub_wire30(4);
	sub_wire1(7, 5)    <= sub_wire30(5);
	sub_wire1(7, 6)    <= sub_wire30(6);
	sub_wire1(7, 7)    <= sub_wire30(7);
	sub_wire1(7, 8)    <= sub_wire30(8);
	sub_wire1(6, 0)    <= sub_wire31(0);
	sub_wire1(6, 1)    <= sub_wire31(1);
	sub_wire1(6, 2)    <= sub_wire31(2);
	sub_wire1(6, 3)    <= sub_wire31(3);
	sub_wire1(6, 4)    <= sub_wire31(4);
	sub_wire1(6, 5)    <= sub_wire31(5);
	sub_wire1(6, 6)    <= sub_wire31(6);
	sub_wire1(6, 7)    <= sub_wire31(7);
	sub_wire1(6, 8)    <= sub_wire31(8);
	sub_wire1(5, 0)    <= sub_wire32(0);
	sub_wire1(5, 1)    <= sub_wire32(1);
	sub_wire1(5, 2)    <= sub_wire32(2);
	sub_wire1(5, 3)    <= sub_wire32(3);
	sub_wire1(5, 4)    <= sub_wire32(4);
	sub_wire1(5, 5)    <= sub_wire32(5);
	sub_wire1(5, 6)    <= sub_wire32(6);
	sub_wire1(5, 7)    <= sub_wire32(7);
	sub_wire1(5, 8)    <= sub_wire32(8);
	sub_wire1(4, 0)    <= sub_wire33(0);
	sub_wire1(4, 1)    <= sub_wire33(1);
	sub_wire1(4, 2)    <= sub_wire33(2);
	sub_wire1(4, 3)    <= sub_wire33(3);
	sub_wire1(4, 4)    <= sub_wire33(4);
	sub_wire1(4, 5)    <= sub_wire33(5);
	sub_wire1(4, 6)    <= sub_wire33(6);
	sub_wire1(4, 7)    <= sub_wire33(7);
	sub_wire1(4, 8)    <= sub_wire33(8);
	sub_wire1(3, 0)    <= sub_wire34(0);
	sub_wire1(3, 1)    <= sub_wire34(1);
	sub_wire1(3, 2)    <= sub_wire34(2);
	sub_wire1(3, 3)    <= sub_wire34(3);
	sub_wire1(3, 4)    <= sub_wire34(4);
	sub_wire1(3, 5)    <= sub_wire34(5);
	sub_wire1(3, 6)    <= sub_wire34(6);
	sub_wire1(3, 7)    <= sub_wire34(7);
	sub_wire1(3, 8)    <= sub_wire34(8);
	sub_wire1(2, 0)    <= sub_wire35(0);
	sub_wire1(2, 1)    <= sub_wire35(1);
	sub_wire1(2, 2)    <= sub_wire35(2);
	sub_wire1(2, 3)    <= sub_wire35(3);
	sub_wire1(2, 4)    <= sub_wire35(4);
	sub_wire1(2, 5)    <= sub_wire35(5);
	sub_wire1(2, 6)    <= sub_wire35(6);
	sub_wire1(2, 7)    <= sub_wire35(7);
	sub_wire1(2, 8)    <= sub_wire35(8);
	sub_wire1(1, 0)    <= sub_wire36(0);
	sub_wire1(1, 1)    <= sub_wire36(1);
	sub_wire1(1, 2)    <= sub_wire36(2);
	sub_wire1(1, 3)    <= sub_wire36(3);
	sub_wire1(1, 4)    <= sub_wire36(4);
	sub_wire1(1, 5)    <= sub_wire36(5);
	sub_wire1(1, 6)    <= sub_wire36(6);
	sub_wire1(1, 7)    <= sub_wire36(7);
	sub_wire1(1, 8)    <= sub_wire36(8);
	sub_wire1(0, 0)    <= sub_wire37(0);
	sub_wire1(0, 1)    <= sub_wire37(1);
	sub_wire1(0, 2)    <= sub_wire37(2);
	sub_wire1(0, 3)    <= sub_wire37(3);
	sub_wire1(0, 4)    <= sub_wire37(4);
	sub_wire1(0, 5)    <= sub_wire37(5);
	sub_wire1(0, 6)    <= sub_wire37(6);
	sub_wire1(0, 7)    <= sub_wire37(7);
	sub_wire1(0, 8)    <= sub_wire37(8);
	result    <= sub_wire38(14 DOWNTO 0);

	parallel_add_component : parallel_add
	GENERIC MAP (
		msw_subtract => "NO",
		pipeline => 1,
		representation => "SIGNED",
		result_alignment => "LSB",
		shift => 0,
		size => 37,
		width => 9,
		widthr => 15,
		lpm_type => "parallel_add"
	)
	PORT MAP (
		aclr => aclr,
		clock => clock,
		data => sub_wire1,
		result => sub_wire38
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: MSW_SUBTRACT STRING "NO"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "1"
-- Retrieval info: CONSTANT: REPRESENTATION STRING "SIGNED"
-- Retrieval info: CONSTANT: RESULT_ALIGNMENT STRING "LSB"
-- Retrieval info: CONSTANT: SHIFT NUMERIC "0"
-- Retrieval info: CONSTANT: SIZE NUMERIC "37"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "9"
-- Retrieval info: CONSTANT: WIDTHR NUMERIC "15"
-- Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT GND "aclr"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT GND "clock"
-- Retrieval info: USED_PORT: data0x 0 0 9 0 INPUT NODEFVAL "data0x[8..0]"
-- Retrieval info: USED_PORT: data10x 0 0 9 0 INPUT NODEFVAL "data10x[8..0]"
-- Retrieval info: USED_PORT: data11x 0 0 9 0 INPUT NODEFVAL "data11x[8..0]"
-- Retrieval info: USED_PORT: data12x 0 0 9 0 INPUT NODEFVAL "data12x[8..0]"
-- Retrieval info: USED_PORT: data13x 0 0 9 0 INPUT NODEFVAL "data13x[8..0]"
-- Retrieval info: USED_PORT: data14x 0 0 9 0 INPUT NODEFVAL "data14x[8..0]"
-- Retrieval info: USED_PORT: data15x 0 0 9 0 INPUT NODEFVAL "data15x[8..0]"
-- Retrieval info: USED_PORT: data16x 0 0 9 0 INPUT NODEFVAL "data16x[8..0]"
-- Retrieval info: USED_PORT: data17x 0 0 9 0 INPUT NODEFVAL "data17x[8..0]"
-- Retrieval info: USED_PORT: data18x 0 0 9 0 INPUT NODEFVAL "data18x[8..0]"
-- Retrieval info: USED_PORT: data19x 0 0 9 0 INPUT NODEFVAL "data19x[8..0]"
-- Retrieval info: USED_PORT: data1x 0 0 9 0 INPUT NODEFVAL "data1x[8..0]"
-- Retrieval info: USED_PORT: data20x 0 0 9 0 INPUT NODEFVAL "data20x[8..0]"
-- Retrieval info: USED_PORT: data21x 0 0 9 0 INPUT NODEFVAL "data21x[8..0]"
-- Retrieval info: USED_PORT: data22x 0 0 9 0 INPUT NODEFVAL "data22x[8..0]"
-- Retrieval info: USED_PORT: data23x 0 0 9 0 INPUT NODEFVAL "data23x[8..0]"
-- Retrieval info: USED_PORT: data24x 0 0 9 0 INPUT NODEFVAL "data24x[8..0]"
-- Retrieval info: USED_PORT: data25x 0 0 9 0 INPUT NODEFVAL "data25x[8..0]"
-- Retrieval info: USED_PORT: data26x 0 0 9 0 INPUT NODEFVAL "data26x[8..0]"
-- Retrieval info: USED_PORT: data27x 0 0 9 0 INPUT NODEFVAL "data27x[8..0]"
-- Retrieval info: USED_PORT: data28x 0 0 9 0 INPUT NODEFVAL "data28x[8..0]"
-- Retrieval info: USED_PORT: data29x 0 0 9 0 INPUT NODEFVAL "data29x[8..0]"
-- Retrieval info: USED_PORT: data2x 0 0 9 0 INPUT NODEFVAL "data2x[8..0]"
-- Retrieval info: USED_PORT: data30x 0 0 9 0 INPUT NODEFVAL "data30x[8..0]"
-- Retrieval info: USED_PORT: data31x 0 0 9 0 INPUT NODEFVAL "data31x[8..0]"
-- Retrieval info: USED_PORT: data32x 0 0 9 0 INPUT NODEFVAL "data32x[8..0]"
-- Retrieval info: USED_PORT: data33x 0 0 9 0 INPUT NODEFVAL "data33x[8..0]"
-- Retrieval info: USED_PORT: data34x 0 0 9 0 INPUT NODEFVAL "data34x[8..0]"
-- Retrieval info: USED_PORT: data35x 0 0 9 0 INPUT NODEFVAL "data35x[8..0]"
-- Retrieval info: USED_PORT: data36x 0 0 9 0 INPUT NODEFVAL "data36x[8..0]"
-- Retrieval info: USED_PORT: data3x 0 0 9 0 INPUT NODEFVAL "data3x[8..0]"
-- Retrieval info: USED_PORT: data4x 0 0 9 0 INPUT NODEFVAL "data4x[8..0]"
-- Retrieval info: USED_PORT: data5x 0 0 9 0 INPUT NODEFVAL "data5x[8..0]"
-- Retrieval info: USED_PORT: data6x 0 0 9 0 INPUT NODEFVAL "data6x[8..0]"
-- Retrieval info: USED_PORT: data7x 0 0 9 0 INPUT NODEFVAL "data7x[8..0]"
-- Retrieval info: USED_PORT: data8x 0 0 9 0 INPUT NODEFVAL "data8x[8..0]"
-- Retrieval info: USED_PORT: data9x 0 0 9 0 INPUT NODEFVAL "data9x[8..0]"
-- Retrieval info: USED_PORT: result 0 0 15 0 OUTPUT NODEFVAL "result[14..0]"
-- Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data 1 0 9 0 data0x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 10 9 0 data10x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 11 9 0 data11x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 12 9 0 data12x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 13 9 0 data13x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 14 9 0 data14x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 15 9 0 data15x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 16 9 0 data16x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 17 9 0 data17x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 18 9 0 data18x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 19 9 0 data19x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 1 9 0 data1x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 20 9 0 data20x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 21 9 0 data21x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 22 9 0 data22x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 23 9 0 data23x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 24 9 0 data24x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 25 9 0 data25x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 26 9 0 data26x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 27 9 0 data27x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 28 9 0 data28x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 29 9 0 data29x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 2 9 0 data2x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 30 9 0 data30x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 31 9 0 data31x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 32 9 0 data32x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 33 9 0 data33x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 34 9 0 data34x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 35 9 0 data35x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 36 9 0 data36x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 3 9 0 data3x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 4 9 0 data4x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 5 9 0 data5x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 6 9 0 data6x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 7 9 0 data7x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 8 9 0 data8x 0 0 9 0
-- Retrieval info: CONNECT: @data 1 9 9 0 data9x 0 0 9 0
-- Retrieval info: CONNECT: result 0 0 15 0 @result 0 0 15 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL Turn_Adder.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Turn_Adder.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Turn_Adder.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Turn_Adder.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Turn_Adder_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
