-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_MUX 

-- ============================================================
-- File Name: MUX8_256b.vhd
-- Megafunction Name(s):
-- 			LPM_MUX
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 15.0.0 Build 145 04/22/2015 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus II License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY MUX8_256b IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data0x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (255 DOWNTO 0)
	);
END MUX8_256b;


ARCHITECTURE SYN OF mux8_256b IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_2D (7 DOWNTO 0, 255 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (255 DOWNTO 0);

BEGIN
	sub_wire8    <= data0x(255 DOWNTO 0);
	sub_wire7    <= data1x(255 DOWNTO 0);
	sub_wire6    <= data2x(255 DOWNTO 0);
	sub_wire5    <= data3x(255 DOWNTO 0);
	sub_wire4    <= data4x(255 DOWNTO 0);
	sub_wire3    <= data5x(255 DOWNTO 0);
	sub_wire2    <= data6x(255 DOWNTO 0);
	sub_wire0    <= data7x(255 DOWNTO 0);
	sub_wire1(7, 0)    <= sub_wire0(0);
	sub_wire1(7, 1)    <= sub_wire0(1);
	sub_wire1(7, 2)    <= sub_wire0(2);
	sub_wire1(7, 3)    <= sub_wire0(3);
	sub_wire1(7, 4)    <= sub_wire0(4);
	sub_wire1(7, 5)    <= sub_wire0(5);
	sub_wire1(7, 6)    <= sub_wire0(6);
	sub_wire1(7, 7)    <= sub_wire0(7);
	sub_wire1(7, 8)    <= sub_wire0(8);
	sub_wire1(7, 9)    <= sub_wire0(9);
	sub_wire1(7, 10)    <= sub_wire0(10);
	sub_wire1(7, 11)    <= sub_wire0(11);
	sub_wire1(7, 12)    <= sub_wire0(12);
	sub_wire1(7, 13)    <= sub_wire0(13);
	sub_wire1(7, 14)    <= sub_wire0(14);
	sub_wire1(7, 15)    <= sub_wire0(15);
	sub_wire1(7, 16)    <= sub_wire0(16);
	sub_wire1(7, 17)    <= sub_wire0(17);
	sub_wire1(7, 18)    <= sub_wire0(18);
	sub_wire1(7, 19)    <= sub_wire0(19);
	sub_wire1(7, 20)    <= sub_wire0(20);
	sub_wire1(7, 21)    <= sub_wire0(21);
	sub_wire1(7, 22)    <= sub_wire0(22);
	sub_wire1(7, 23)    <= sub_wire0(23);
	sub_wire1(7, 24)    <= sub_wire0(24);
	sub_wire1(7, 25)    <= sub_wire0(25);
	sub_wire1(7, 26)    <= sub_wire0(26);
	sub_wire1(7, 27)    <= sub_wire0(27);
	sub_wire1(7, 28)    <= sub_wire0(28);
	sub_wire1(7, 29)    <= sub_wire0(29);
	sub_wire1(7, 30)    <= sub_wire0(30);
	sub_wire1(7, 31)    <= sub_wire0(31);
	sub_wire1(7, 32)    <= sub_wire0(32);
	sub_wire1(7, 33)    <= sub_wire0(33);
	sub_wire1(7, 34)    <= sub_wire0(34);
	sub_wire1(7, 35)    <= sub_wire0(35);
	sub_wire1(7, 36)    <= sub_wire0(36);
	sub_wire1(7, 37)    <= sub_wire0(37);
	sub_wire1(7, 38)    <= sub_wire0(38);
	sub_wire1(7, 39)    <= sub_wire0(39);
	sub_wire1(7, 40)    <= sub_wire0(40);
	sub_wire1(7, 41)    <= sub_wire0(41);
	sub_wire1(7, 42)    <= sub_wire0(42);
	sub_wire1(7, 43)    <= sub_wire0(43);
	sub_wire1(7, 44)    <= sub_wire0(44);
	sub_wire1(7, 45)    <= sub_wire0(45);
	sub_wire1(7, 46)    <= sub_wire0(46);
	sub_wire1(7, 47)    <= sub_wire0(47);
	sub_wire1(7, 48)    <= sub_wire0(48);
	sub_wire1(7, 49)    <= sub_wire0(49);
	sub_wire1(7, 50)    <= sub_wire0(50);
	sub_wire1(7, 51)    <= sub_wire0(51);
	sub_wire1(7, 52)    <= sub_wire0(52);
	sub_wire1(7, 53)    <= sub_wire0(53);
	sub_wire1(7, 54)    <= sub_wire0(54);
	sub_wire1(7, 55)    <= sub_wire0(55);
	sub_wire1(7, 56)    <= sub_wire0(56);
	sub_wire1(7, 57)    <= sub_wire0(57);
	sub_wire1(7, 58)    <= sub_wire0(58);
	sub_wire1(7, 59)    <= sub_wire0(59);
	sub_wire1(7, 60)    <= sub_wire0(60);
	sub_wire1(7, 61)    <= sub_wire0(61);
	sub_wire1(7, 62)    <= sub_wire0(62);
	sub_wire1(7, 63)    <= sub_wire0(63);
	sub_wire1(7, 64)    <= sub_wire0(64);
	sub_wire1(7, 65)    <= sub_wire0(65);
	sub_wire1(7, 66)    <= sub_wire0(66);
	sub_wire1(7, 67)    <= sub_wire0(67);
	sub_wire1(7, 68)    <= sub_wire0(68);
	sub_wire1(7, 69)    <= sub_wire0(69);
	sub_wire1(7, 70)    <= sub_wire0(70);
	sub_wire1(7, 71)    <= sub_wire0(71);
	sub_wire1(7, 72)    <= sub_wire0(72);
	sub_wire1(7, 73)    <= sub_wire0(73);
	sub_wire1(7, 74)    <= sub_wire0(74);
	sub_wire1(7, 75)    <= sub_wire0(75);
	sub_wire1(7, 76)    <= sub_wire0(76);
	sub_wire1(7, 77)    <= sub_wire0(77);
	sub_wire1(7, 78)    <= sub_wire0(78);
	sub_wire1(7, 79)    <= sub_wire0(79);
	sub_wire1(7, 80)    <= sub_wire0(80);
	sub_wire1(7, 81)    <= sub_wire0(81);
	sub_wire1(7, 82)    <= sub_wire0(82);
	sub_wire1(7, 83)    <= sub_wire0(83);
	sub_wire1(7, 84)    <= sub_wire0(84);
	sub_wire1(7, 85)    <= sub_wire0(85);
	sub_wire1(7, 86)    <= sub_wire0(86);
	sub_wire1(7, 87)    <= sub_wire0(87);
	sub_wire1(7, 88)    <= sub_wire0(88);
	sub_wire1(7, 89)    <= sub_wire0(89);
	sub_wire1(7, 90)    <= sub_wire0(90);
	sub_wire1(7, 91)    <= sub_wire0(91);
	sub_wire1(7, 92)    <= sub_wire0(92);
	sub_wire1(7, 93)    <= sub_wire0(93);
	sub_wire1(7, 94)    <= sub_wire0(94);
	sub_wire1(7, 95)    <= sub_wire0(95);
	sub_wire1(7, 96)    <= sub_wire0(96);
	sub_wire1(7, 97)    <= sub_wire0(97);
	sub_wire1(7, 98)    <= sub_wire0(98);
	sub_wire1(7, 99)    <= sub_wire0(99);
	sub_wire1(7, 100)    <= sub_wire0(100);
	sub_wire1(7, 101)    <= sub_wire0(101);
	sub_wire1(7, 102)    <= sub_wire0(102);
	sub_wire1(7, 103)    <= sub_wire0(103);
	sub_wire1(7, 104)    <= sub_wire0(104);
	sub_wire1(7, 105)    <= sub_wire0(105);
	sub_wire1(7, 106)    <= sub_wire0(106);
	sub_wire1(7, 107)    <= sub_wire0(107);
	sub_wire1(7, 108)    <= sub_wire0(108);
	sub_wire1(7, 109)    <= sub_wire0(109);
	sub_wire1(7, 110)    <= sub_wire0(110);
	sub_wire1(7, 111)    <= sub_wire0(111);
	sub_wire1(7, 112)    <= sub_wire0(112);
	sub_wire1(7, 113)    <= sub_wire0(113);
	sub_wire1(7, 114)    <= sub_wire0(114);
	sub_wire1(7, 115)    <= sub_wire0(115);
	sub_wire1(7, 116)    <= sub_wire0(116);
	sub_wire1(7, 117)    <= sub_wire0(117);
	sub_wire1(7, 118)    <= sub_wire0(118);
	sub_wire1(7, 119)    <= sub_wire0(119);
	sub_wire1(7, 120)    <= sub_wire0(120);
	sub_wire1(7, 121)    <= sub_wire0(121);
	sub_wire1(7, 122)    <= sub_wire0(122);
	sub_wire1(7, 123)    <= sub_wire0(123);
	sub_wire1(7, 124)    <= sub_wire0(124);
	sub_wire1(7, 125)    <= sub_wire0(125);
	sub_wire1(7, 126)    <= sub_wire0(126);
	sub_wire1(7, 127)    <= sub_wire0(127);
	sub_wire1(7, 128)    <= sub_wire0(128);
	sub_wire1(7, 129)    <= sub_wire0(129);
	sub_wire1(7, 130)    <= sub_wire0(130);
	sub_wire1(7, 131)    <= sub_wire0(131);
	sub_wire1(7, 132)    <= sub_wire0(132);
	sub_wire1(7, 133)    <= sub_wire0(133);
	sub_wire1(7, 134)    <= sub_wire0(134);
	sub_wire1(7, 135)    <= sub_wire0(135);
	sub_wire1(7, 136)    <= sub_wire0(136);
	sub_wire1(7, 137)    <= sub_wire0(137);
	sub_wire1(7, 138)    <= sub_wire0(138);
	sub_wire1(7, 139)    <= sub_wire0(139);
	sub_wire1(7, 140)    <= sub_wire0(140);
	sub_wire1(7, 141)    <= sub_wire0(141);
	sub_wire1(7, 142)    <= sub_wire0(142);
	sub_wire1(7, 143)    <= sub_wire0(143);
	sub_wire1(7, 144)    <= sub_wire0(144);
	sub_wire1(7, 145)    <= sub_wire0(145);
	sub_wire1(7, 146)    <= sub_wire0(146);
	sub_wire1(7, 147)    <= sub_wire0(147);
	sub_wire1(7, 148)    <= sub_wire0(148);
	sub_wire1(7, 149)    <= sub_wire0(149);
	sub_wire1(7, 150)    <= sub_wire0(150);
	sub_wire1(7, 151)    <= sub_wire0(151);
	sub_wire1(7, 152)    <= sub_wire0(152);
	sub_wire1(7, 153)    <= sub_wire0(153);
	sub_wire1(7, 154)    <= sub_wire0(154);
	sub_wire1(7, 155)    <= sub_wire0(155);
	sub_wire1(7, 156)    <= sub_wire0(156);
	sub_wire1(7, 157)    <= sub_wire0(157);
	sub_wire1(7, 158)    <= sub_wire0(158);
	sub_wire1(7, 159)    <= sub_wire0(159);
	sub_wire1(7, 160)    <= sub_wire0(160);
	sub_wire1(7, 161)    <= sub_wire0(161);
	sub_wire1(7, 162)    <= sub_wire0(162);
	sub_wire1(7, 163)    <= sub_wire0(163);
	sub_wire1(7, 164)    <= sub_wire0(164);
	sub_wire1(7, 165)    <= sub_wire0(165);
	sub_wire1(7, 166)    <= sub_wire0(166);
	sub_wire1(7, 167)    <= sub_wire0(167);
	sub_wire1(7, 168)    <= sub_wire0(168);
	sub_wire1(7, 169)    <= sub_wire0(169);
	sub_wire1(7, 170)    <= sub_wire0(170);
	sub_wire1(7, 171)    <= sub_wire0(171);
	sub_wire1(7, 172)    <= sub_wire0(172);
	sub_wire1(7, 173)    <= sub_wire0(173);
	sub_wire1(7, 174)    <= sub_wire0(174);
	sub_wire1(7, 175)    <= sub_wire0(175);
	sub_wire1(7, 176)    <= sub_wire0(176);
	sub_wire1(7, 177)    <= sub_wire0(177);
	sub_wire1(7, 178)    <= sub_wire0(178);
	sub_wire1(7, 179)    <= sub_wire0(179);
	sub_wire1(7, 180)    <= sub_wire0(180);
	sub_wire1(7, 181)    <= sub_wire0(181);
	sub_wire1(7, 182)    <= sub_wire0(182);
	sub_wire1(7, 183)    <= sub_wire0(183);
	sub_wire1(7, 184)    <= sub_wire0(184);
	sub_wire1(7, 185)    <= sub_wire0(185);
	sub_wire1(7, 186)    <= sub_wire0(186);
	sub_wire1(7, 187)    <= sub_wire0(187);
	sub_wire1(7, 188)    <= sub_wire0(188);
	sub_wire1(7, 189)    <= sub_wire0(189);
	sub_wire1(7, 190)    <= sub_wire0(190);
	sub_wire1(7, 191)    <= sub_wire0(191);
	sub_wire1(7, 192)    <= sub_wire0(192);
	sub_wire1(7, 193)    <= sub_wire0(193);
	sub_wire1(7, 194)    <= sub_wire0(194);
	sub_wire1(7, 195)    <= sub_wire0(195);
	sub_wire1(7, 196)    <= sub_wire0(196);
	sub_wire1(7, 197)    <= sub_wire0(197);
	sub_wire1(7, 198)    <= sub_wire0(198);
	sub_wire1(7, 199)    <= sub_wire0(199);
	sub_wire1(7, 200)    <= sub_wire0(200);
	sub_wire1(7, 201)    <= sub_wire0(201);
	sub_wire1(7, 202)    <= sub_wire0(202);
	sub_wire1(7, 203)    <= sub_wire0(203);
	sub_wire1(7, 204)    <= sub_wire0(204);
	sub_wire1(7, 205)    <= sub_wire0(205);
	sub_wire1(7, 206)    <= sub_wire0(206);
	sub_wire1(7, 207)    <= sub_wire0(207);
	sub_wire1(7, 208)    <= sub_wire0(208);
	sub_wire1(7, 209)    <= sub_wire0(209);
	sub_wire1(7, 210)    <= sub_wire0(210);
	sub_wire1(7, 211)    <= sub_wire0(211);
	sub_wire1(7, 212)    <= sub_wire0(212);
	sub_wire1(7, 213)    <= sub_wire0(213);
	sub_wire1(7, 214)    <= sub_wire0(214);
	sub_wire1(7, 215)    <= sub_wire0(215);
	sub_wire1(7, 216)    <= sub_wire0(216);
	sub_wire1(7, 217)    <= sub_wire0(217);
	sub_wire1(7, 218)    <= sub_wire0(218);
	sub_wire1(7, 219)    <= sub_wire0(219);
	sub_wire1(7, 220)    <= sub_wire0(220);
	sub_wire1(7, 221)    <= sub_wire0(221);
	sub_wire1(7, 222)    <= sub_wire0(222);
	sub_wire1(7, 223)    <= sub_wire0(223);
	sub_wire1(7, 224)    <= sub_wire0(224);
	sub_wire1(7, 225)    <= sub_wire0(225);
	sub_wire1(7, 226)    <= sub_wire0(226);
	sub_wire1(7, 227)    <= sub_wire0(227);
	sub_wire1(7, 228)    <= sub_wire0(228);
	sub_wire1(7, 229)    <= sub_wire0(229);
	sub_wire1(7, 230)    <= sub_wire0(230);
	sub_wire1(7, 231)    <= sub_wire0(231);
	sub_wire1(7, 232)    <= sub_wire0(232);
	sub_wire1(7, 233)    <= sub_wire0(233);
	sub_wire1(7, 234)    <= sub_wire0(234);
	sub_wire1(7, 235)    <= sub_wire0(235);
	sub_wire1(7, 236)    <= sub_wire0(236);
	sub_wire1(7, 237)    <= sub_wire0(237);
	sub_wire1(7, 238)    <= sub_wire0(238);
	sub_wire1(7, 239)    <= sub_wire0(239);
	sub_wire1(7, 240)    <= sub_wire0(240);
	sub_wire1(7, 241)    <= sub_wire0(241);
	sub_wire1(7, 242)    <= sub_wire0(242);
	sub_wire1(7, 243)    <= sub_wire0(243);
	sub_wire1(7, 244)    <= sub_wire0(244);
	sub_wire1(7, 245)    <= sub_wire0(245);
	sub_wire1(7, 246)    <= sub_wire0(246);
	sub_wire1(7, 247)    <= sub_wire0(247);
	sub_wire1(7, 248)    <= sub_wire0(248);
	sub_wire1(7, 249)    <= sub_wire0(249);
	sub_wire1(7, 250)    <= sub_wire0(250);
	sub_wire1(7, 251)    <= sub_wire0(251);
	sub_wire1(7, 252)    <= sub_wire0(252);
	sub_wire1(7, 253)    <= sub_wire0(253);
	sub_wire1(7, 254)    <= sub_wire0(254);
	sub_wire1(7, 255)    <= sub_wire0(255);
	sub_wire1(6, 0)    <= sub_wire2(0);
	sub_wire1(6, 1)    <= sub_wire2(1);
	sub_wire1(6, 2)    <= sub_wire2(2);
	sub_wire1(6, 3)    <= sub_wire2(3);
	sub_wire1(6, 4)    <= sub_wire2(4);
	sub_wire1(6, 5)    <= sub_wire2(5);
	sub_wire1(6, 6)    <= sub_wire2(6);
	sub_wire1(6, 7)    <= sub_wire2(7);
	sub_wire1(6, 8)    <= sub_wire2(8);
	sub_wire1(6, 9)    <= sub_wire2(9);
	sub_wire1(6, 10)    <= sub_wire2(10);
	sub_wire1(6, 11)    <= sub_wire2(11);
	sub_wire1(6, 12)    <= sub_wire2(12);
	sub_wire1(6, 13)    <= sub_wire2(13);
	sub_wire1(6, 14)    <= sub_wire2(14);
	sub_wire1(6, 15)    <= sub_wire2(15);
	sub_wire1(6, 16)    <= sub_wire2(16);
	sub_wire1(6, 17)    <= sub_wire2(17);
	sub_wire1(6, 18)    <= sub_wire2(18);
	sub_wire1(6, 19)    <= sub_wire2(19);
	sub_wire1(6, 20)    <= sub_wire2(20);
	sub_wire1(6, 21)    <= sub_wire2(21);
	sub_wire1(6, 22)    <= sub_wire2(22);
	sub_wire1(6, 23)    <= sub_wire2(23);
	sub_wire1(6, 24)    <= sub_wire2(24);
	sub_wire1(6, 25)    <= sub_wire2(25);
	sub_wire1(6, 26)    <= sub_wire2(26);
	sub_wire1(6, 27)    <= sub_wire2(27);
	sub_wire1(6, 28)    <= sub_wire2(28);
	sub_wire1(6, 29)    <= sub_wire2(29);
	sub_wire1(6, 30)    <= sub_wire2(30);
	sub_wire1(6, 31)    <= sub_wire2(31);
	sub_wire1(6, 32)    <= sub_wire2(32);
	sub_wire1(6, 33)    <= sub_wire2(33);
	sub_wire1(6, 34)    <= sub_wire2(34);
	sub_wire1(6, 35)    <= sub_wire2(35);
	sub_wire1(6, 36)    <= sub_wire2(36);
	sub_wire1(6, 37)    <= sub_wire2(37);
	sub_wire1(6, 38)    <= sub_wire2(38);
	sub_wire1(6, 39)    <= sub_wire2(39);
	sub_wire1(6, 40)    <= sub_wire2(40);
	sub_wire1(6, 41)    <= sub_wire2(41);
	sub_wire1(6, 42)    <= sub_wire2(42);
	sub_wire1(6, 43)    <= sub_wire2(43);
	sub_wire1(6, 44)    <= sub_wire2(44);
	sub_wire1(6, 45)    <= sub_wire2(45);
	sub_wire1(6, 46)    <= sub_wire2(46);
	sub_wire1(6, 47)    <= sub_wire2(47);
	sub_wire1(6, 48)    <= sub_wire2(48);
	sub_wire1(6, 49)    <= sub_wire2(49);
	sub_wire1(6, 50)    <= sub_wire2(50);
	sub_wire1(6, 51)    <= sub_wire2(51);
	sub_wire1(6, 52)    <= sub_wire2(52);
	sub_wire1(6, 53)    <= sub_wire2(53);
	sub_wire1(6, 54)    <= sub_wire2(54);
	sub_wire1(6, 55)    <= sub_wire2(55);
	sub_wire1(6, 56)    <= sub_wire2(56);
	sub_wire1(6, 57)    <= sub_wire2(57);
	sub_wire1(6, 58)    <= sub_wire2(58);
	sub_wire1(6, 59)    <= sub_wire2(59);
	sub_wire1(6, 60)    <= sub_wire2(60);
	sub_wire1(6, 61)    <= sub_wire2(61);
	sub_wire1(6, 62)    <= sub_wire2(62);
	sub_wire1(6, 63)    <= sub_wire2(63);
	sub_wire1(6, 64)    <= sub_wire2(64);
	sub_wire1(6, 65)    <= sub_wire2(65);
	sub_wire1(6, 66)    <= sub_wire2(66);
	sub_wire1(6, 67)    <= sub_wire2(67);
	sub_wire1(6, 68)    <= sub_wire2(68);
	sub_wire1(6, 69)    <= sub_wire2(69);
	sub_wire1(6, 70)    <= sub_wire2(70);
	sub_wire1(6, 71)    <= sub_wire2(71);
	sub_wire1(6, 72)    <= sub_wire2(72);
	sub_wire1(6, 73)    <= sub_wire2(73);
	sub_wire1(6, 74)    <= sub_wire2(74);
	sub_wire1(6, 75)    <= sub_wire2(75);
	sub_wire1(6, 76)    <= sub_wire2(76);
	sub_wire1(6, 77)    <= sub_wire2(77);
	sub_wire1(6, 78)    <= sub_wire2(78);
	sub_wire1(6, 79)    <= sub_wire2(79);
	sub_wire1(6, 80)    <= sub_wire2(80);
	sub_wire1(6, 81)    <= sub_wire2(81);
	sub_wire1(6, 82)    <= sub_wire2(82);
	sub_wire1(6, 83)    <= sub_wire2(83);
	sub_wire1(6, 84)    <= sub_wire2(84);
	sub_wire1(6, 85)    <= sub_wire2(85);
	sub_wire1(6, 86)    <= sub_wire2(86);
	sub_wire1(6, 87)    <= sub_wire2(87);
	sub_wire1(6, 88)    <= sub_wire2(88);
	sub_wire1(6, 89)    <= sub_wire2(89);
	sub_wire1(6, 90)    <= sub_wire2(90);
	sub_wire1(6, 91)    <= sub_wire2(91);
	sub_wire1(6, 92)    <= sub_wire2(92);
	sub_wire1(6, 93)    <= sub_wire2(93);
	sub_wire1(6, 94)    <= sub_wire2(94);
	sub_wire1(6, 95)    <= sub_wire2(95);
	sub_wire1(6, 96)    <= sub_wire2(96);
	sub_wire1(6, 97)    <= sub_wire2(97);
	sub_wire1(6, 98)    <= sub_wire2(98);
	sub_wire1(6, 99)    <= sub_wire2(99);
	sub_wire1(6, 100)    <= sub_wire2(100);
	sub_wire1(6, 101)    <= sub_wire2(101);
	sub_wire1(6, 102)    <= sub_wire2(102);
	sub_wire1(6, 103)    <= sub_wire2(103);
	sub_wire1(6, 104)    <= sub_wire2(104);
	sub_wire1(6, 105)    <= sub_wire2(105);
	sub_wire1(6, 106)    <= sub_wire2(106);
	sub_wire1(6, 107)    <= sub_wire2(107);
	sub_wire1(6, 108)    <= sub_wire2(108);
	sub_wire1(6, 109)    <= sub_wire2(109);
	sub_wire1(6, 110)    <= sub_wire2(110);
	sub_wire1(6, 111)    <= sub_wire2(111);
	sub_wire1(6, 112)    <= sub_wire2(112);
	sub_wire1(6, 113)    <= sub_wire2(113);
	sub_wire1(6, 114)    <= sub_wire2(114);
	sub_wire1(6, 115)    <= sub_wire2(115);
	sub_wire1(6, 116)    <= sub_wire2(116);
	sub_wire1(6, 117)    <= sub_wire2(117);
	sub_wire1(6, 118)    <= sub_wire2(118);
	sub_wire1(6, 119)    <= sub_wire2(119);
	sub_wire1(6, 120)    <= sub_wire2(120);
	sub_wire1(6, 121)    <= sub_wire2(121);
	sub_wire1(6, 122)    <= sub_wire2(122);
	sub_wire1(6, 123)    <= sub_wire2(123);
	sub_wire1(6, 124)    <= sub_wire2(124);
	sub_wire1(6, 125)    <= sub_wire2(125);
	sub_wire1(6, 126)    <= sub_wire2(126);
	sub_wire1(6, 127)    <= sub_wire2(127);
	sub_wire1(6, 128)    <= sub_wire2(128);
	sub_wire1(6, 129)    <= sub_wire2(129);
	sub_wire1(6, 130)    <= sub_wire2(130);
	sub_wire1(6, 131)    <= sub_wire2(131);
	sub_wire1(6, 132)    <= sub_wire2(132);
	sub_wire1(6, 133)    <= sub_wire2(133);
	sub_wire1(6, 134)    <= sub_wire2(134);
	sub_wire1(6, 135)    <= sub_wire2(135);
	sub_wire1(6, 136)    <= sub_wire2(136);
	sub_wire1(6, 137)    <= sub_wire2(137);
	sub_wire1(6, 138)    <= sub_wire2(138);
	sub_wire1(6, 139)    <= sub_wire2(139);
	sub_wire1(6, 140)    <= sub_wire2(140);
	sub_wire1(6, 141)    <= sub_wire2(141);
	sub_wire1(6, 142)    <= sub_wire2(142);
	sub_wire1(6, 143)    <= sub_wire2(143);
	sub_wire1(6, 144)    <= sub_wire2(144);
	sub_wire1(6, 145)    <= sub_wire2(145);
	sub_wire1(6, 146)    <= sub_wire2(146);
	sub_wire1(6, 147)    <= sub_wire2(147);
	sub_wire1(6, 148)    <= sub_wire2(148);
	sub_wire1(6, 149)    <= sub_wire2(149);
	sub_wire1(6, 150)    <= sub_wire2(150);
	sub_wire1(6, 151)    <= sub_wire2(151);
	sub_wire1(6, 152)    <= sub_wire2(152);
	sub_wire1(6, 153)    <= sub_wire2(153);
	sub_wire1(6, 154)    <= sub_wire2(154);
	sub_wire1(6, 155)    <= sub_wire2(155);
	sub_wire1(6, 156)    <= sub_wire2(156);
	sub_wire1(6, 157)    <= sub_wire2(157);
	sub_wire1(6, 158)    <= sub_wire2(158);
	sub_wire1(6, 159)    <= sub_wire2(159);
	sub_wire1(6, 160)    <= sub_wire2(160);
	sub_wire1(6, 161)    <= sub_wire2(161);
	sub_wire1(6, 162)    <= sub_wire2(162);
	sub_wire1(6, 163)    <= sub_wire2(163);
	sub_wire1(6, 164)    <= sub_wire2(164);
	sub_wire1(6, 165)    <= sub_wire2(165);
	sub_wire1(6, 166)    <= sub_wire2(166);
	sub_wire1(6, 167)    <= sub_wire2(167);
	sub_wire1(6, 168)    <= sub_wire2(168);
	sub_wire1(6, 169)    <= sub_wire2(169);
	sub_wire1(6, 170)    <= sub_wire2(170);
	sub_wire1(6, 171)    <= sub_wire2(171);
	sub_wire1(6, 172)    <= sub_wire2(172);
	sub_wire1(6, 173)    <= sub_wire2(173);
	sub_wire1(6, 174)    <= sub_wire2(174);
	sub_wire1(6, 175)    <= sub_wire2(175);
	sub_wire1(6, 176)    <= sub_wire2(176);
	sub_wire1(6, 177)    <= sub_wire2(177);
	sub_wire1(6, 178)    <= sub_wire2(178);
	sub_wire1(6, 179)    <= sub_wire2(179);
	sub_wire1(6, 180)    <= sub_wire2(180);
	sub_wire1(6, 181)    <= sub_wire2(181);
	sub_wire1(6, 182)    <= sub_wire2(182);
	sub_wire1(6, 183)    <= sub_wire2(183);
	sub_wire1(6, 184)    <= sub_wire2(184);
	sub_wire1(6, 185)    <= sub_wire2(185);
	sub_wire1(6, 186)    <= sub_wire2(186);
	sub_wire1(6, 187)    <= sub_wire2(187);
	sub_wire1(6, 188)    <= sub_wire2(188);
	sub_wire1(6, 189)    <= sub_wire2(189);
	sub_wire1(6, 190)    <= sub_wire2(190);
	sub_wire1(6, 191)    <= sub_wire2(191);
	sub_wire1(6, 192)    <= sub_wire2(192);
	sub_wire1(6, 193)    <= sub_wire2(193);
	sub_wire1(6, 194)    <= sub_wire2(194);
	sub_wire1(6, 195)    <= sub_wire2(195);
	sub_wire1(6, 196)    <= sub_wire2(196);
	sub_wire1(6, 197)    <= sub_wire2(197);
	sub_wire1(6, 198)    <= sub_wire2(198);
	sub_wire1(6, 199)    <= sub_wire2(199);
	sub_wire1(6, 200)    <= sub_wire2(200);
	sub_wire1(6, 201)    <= sub_wire2(201);
	sub_wire1(6, 202)    <= sub_wire2(202);
	sub_wire1(6, 203)    <= sub_wire2(203);
	sub_wire1(6, 204)    <= sub_wire2(204);
	sub_wire1(6, 205)    <= sub_wire2(205);
	sub_wire1(6, 206)    <= sub_wire2(206);
	sub_wire1(6, 207)    <= sub_wire2(207);
	sub_wire1(6, 208)    <= sub_wire2(208);
	sub_wire1(6, 209)    <= sub_wire2(209);
	sub_wire1(6, 210)    <= sub_wire2(210);
	sub_wire1(6, 211)    <= sub_wire2(211);
	sub_wire1(6, 212)    <= sub_wire2(212);
	sub_wire1(6, 213)    <= sub_wire2(213);
	sub_wire1(6, 214)    <= sub_wire2(214);
	sub_wire1(6, 215)    <= sub_wire2(215);
	sub_wire1(6, 216)    <= sub_wire2(216);
	sub_wire1(6, 217)    <= sub_wire2(217);
	sub_wire1(6, 218)    <= sub_wire2(218);
	sub_wire1(6, 219)    <= sub_wire2(219);
	sub_wire1(6, 220)    <= sub_wire2(220);
	sub_wire1(6, 221)    <= sub_wire2(221);
	sub_wire1(6, 222)    <= sub_wire2(222);
	sub_wire1(6, 223)    <= sub_wire2(223);
	sub_wire1(6, 224)    <= sub_wire2(224);
	sub_wire1(6, 225)    <= sub_wire2(225);
	sub_wire1(6, 226)    <= sub_wire2(226);
	sub_wire1(6, 227)    <= sub_wire2(227);
	sub_wire1(6, 228)    <= sub_wire2(228);
	sub_wire1(6, 229)    <= sub_wire2(229);
	sub_wire1(6, 230)    <= sub_wire2(230);
	sub_wire1(6, 231)    <= sub_wire2(231);
	sub_wire1(6, 232)    <= sub_wire2(232);
	sub_wire1(6, 233)    <= sub_wire2(233);
	sub_wire1(6, 234)    <= sub_wire2(234);
	sub_wire1(6, 235)    <= sub_wire2(235);
	sub_wire1(6, 236)    <= sub_wire2(236);
	sub_wire1(6, 237)    <= sub_wire2(237);
	sub_wire1(6, 238)    <= sub_wire2(238);
	sub_wire1(6, 239)    <= sub_wire2(239);
	sub_wire1(6, 240)    <= sub_wire2(240);
	sub_wire1(6, 241)    <= sub_wire2(241);
	sub_wire1(6, 242)    <= sub_wire2(242);
	sub_wire1(6, 243)    <= sub_wire2(243);
	sub_wire1(6, 244)    <= sub_wire2(244);
	sub_wire1(6, 245)    <= sub_wire2(245);
	sub_wire1(6, 246)    <= sub_wire2(246);
	sub_wire1(6, 247)    <= sub_wire2(247);
	sub_wire1(6, 248)    <= sub_wire2(248);
	sub_wire1(6, 249)    <= sub_wire2(249);
	sub_wire1(6, 250)    <= sub_wire2(250);
	sub_wire1(6, 251)    <= sub_wire2(251);
	sub_wire1(6, 252)    <= sub_wire2(252);
	sub_wire1(6, 253)    <= sub_wire2(253);
	sub_wire1(6, 254)    <= sub_wire2(254);
	sub_wire1(6, 255)    <= sub_wire2(255);
	sub_wire1(5, 0)    <= sub_wire3(0);
	sub_wire1(5, 1)    <= sub_wire3(1);
	sub_wire1(5, 2)    <= sub_wire3(2);
	sub_wire1(5, 3)    <= sub_wire3(3);
	sub_wire1(5, 4)    <= sub_wire3(4);
	sub_wire1(5, 5)    <= sub_wire3(5);
	sub_wire1(5, 6)    <= sub_wire3(6);
	sub_wire1(5, 7)    <= sub_wire3(7);
	sub_wire1(5, 8)    <= sub_wire3(8);
	sub_wire1(5, 9)    <= sub_wire3(9);
	sub_wire1(5, 10)    <= sub_wire3(10);
	sub_wire1(5, 11)    <= sub_wire3(11);
	sub_wire1(5, 12)    <= sub_wire3(12);
	sub_wire1(5, 13)    <= sub_wire3(13);
	sub_wire1(5, 14)    <= sub_wire3(14);
	sub_wire1(5, 15)    <= sub_wire3(15);
	sub_wire1(5, 16)    <= sub_wire3(16);
	sub_wire1(5, 17)    <= sub_wire3(17);
	sub_wire1(5, 18)    <= sub_wire3(18);
	sub_wire1(5, 19)    <= sub_wire3(19);
	sub_wire1(5, 20)    <= sub_wire3(20);
	sub_wire1(5, 21)    <= sub_wire3(21);
	sub_wire1(5, 22)    <= sub_wire3(22);
	sub_wire1(5, 23)    <= sub_wire3(23);
	sub_wire1(5, 24)    <= sub_wire3(24);
	sub_wire1(5, 25)    <= sub_wire3(25);
	sub_wire1(5, 26)    <= sub_wire3(26);
	sub_wire1(5, 27)    <= sub_wire3(27);
	sub_wire1(5, 28)    <= sub_wire3(28);
	sub_wire1(5, 29)    <= sub_wire3(29);
	sub_wire1(5, 30)    <= sub_wire3(30);
	sub_wire1(5, 31)    <= sub_wire3(31);
	sub_wire1(5, 32)    <= sub_wire3(32);
	sub_wire1(5, 33)    <= sub_wire3(33);
	sub_wire1(5, 34)    <= sub_wire3(34);
	sub_wire1(5, 35)    <= sub_wire3(35);
	sub_wire1(5, 36)    <= sub_wire3(36);
	sub_wire1(5, 37)    <= sub_wire3(37);
	sub_wire1(5, 38)    <= sub_wire3(38);
	sub_wire1(5, 39)    <= sub_wire3(39);
	sub_wire1(5, 40)    <= sub_wire3(40);
	sub_wire1(5, 41)    <= sub_wire3(41);
	sub_wire1(5, 42)    <= sub_wire3(42);
	sub_wire1(5, 43)    <= sub_wire3(43);
	sub_wire1(5, 44)    <= sub_wire3(44);
	sub_wire1(5, 45)    <= sub_wire3(45);
	sub_wire1(5, 46)    <= sub_wire3(46);
	sub_wire1(5, 47)    <= sub_wire3(47);
	sub_wire1(5, 48)    <= sub_wire3(48);
	sub_wire1(5, 49)    <= sub_wire3(49);
	sub_wire1(5, 50)    <= sub_wire3(50);
	sub_wire1(5, 51)    <= sub_wire3(51);
	sub_wire1(5, 52)    <= sub_wire3(52);
	sub_wire1(5, 53)    <= sub_wire3(53);
	sub_wire1(5, 54)    <= sub_wire3(54);
	sub_wire1(5, 55)    <= sub_wire3(55);
	sub_wire1(5, 56)    <= sub_wire3(56);
	sub_wire1(5, 57)    <= sub_wire3(57);
	sub_wire1(5, 58)    <= sub_wire3(58);
	sub_wire1(5, 59)    <= sub_wire3(59);
	sub_wire1(5, 60)    <= sub_wire3(60);
	sub_wire1(5, 61)    <= sub_wire3(61);
	sub_wire1(5, 62)    <= sub_wire3(62);
	sub_wire1(5, 63)    <= sub_wire3(63);
	sub_wire1(5, 64)    <= sub_wire3(64);
	sub_wire1(5, 65)    <= sub_wire3(65);
	sub_wire1(5, 66)    <= sub_wire3(66);
	sub_wire1(5, 67)    <= sub_wire3(67);
	sub_wire1(5, 68)    <= sub_wire3(68);
	sub_wire1(5, 69)    <= sub_wire3(69);
	sub_wire1(5, 70)    <= sub_wire3(70);
	sub_wire1(5, 71)    <= sub_wire3(71);
	sub_wire1(5, 72)    <= sub_wire3(72);
	sub_wire1(5, 73)    <= sub_wire3(73);
	sub_wire1(5, 74)    <= sub_wire3(74);
	sub_wire1(5, 75)    <= sub_wire3(75);
	sub_wire1(5, 76)    <= sub_wire3(76);
	sub_wire1(5, 77)    <= sub_wire3(77);
	sub_wire1(5, 78)    <= sub_wire3(78);
	sub_wire1(5, 79)    <= sub_wire3(79);
	sub_wire1(5, 80)    <= sub_wire3(80);
	sub_wire1(5, 81)    <= sub_wire3(81);
	sub_wire1(5, 82)    <= sub_wire3(82);
	sub_wire1(5, 83)    <= sub_wire3(83);
	sub_wire1(5, 84)    <= sub_wire3(84);
	sub_wire1(5, 85)    <= sub_wire3(85);
	sub_wire1(5, 86)    <= sub_wire3(86);
	sub_wire1(5, 87)    <= sub_wire3(87);
	sub_wire1(5, 88)    <= sub_wire3(88);
	sub_wire1(5, 89)    <= sub_wire3(89);
	sub_wire1(5, 90)    <= sub_wire3(90);
	sub_wire1(5, 91)    <= sub_wire3(91);
	sub_wire1(5, 92)    <= sub_wire3(92);
	sub_wire1(5, 93)    <= sub_wire3(93);
	sub_wire1(5, 94)    <= sub_wire3(94);
	sub_wire1(5, 95)    <= sub_wire3(95);
	sub_wire1(5, 96)    <= sub_wire3(96);
	sub_wire1(5, 97)    <= sub_wire3(97);
	sub_wire1(5, 98)    <= sub_wire3(98);
	sub_wire1(5, 99)    <= sub_wire3(99);
	sub_wire1(5, 100)    <= sub_wire3(100);
	sub_wire1(5, 101)    <= sub_wire3(101);
	sub_wire1(5, 102)    <= sub_wire3(102);
	sub_wire1(5, 103)    <= sub_wire3(103);
	sub_wire1(5, 104)    <= sub_wire3(104);
	sub_wire1(5, 105)    <= sub_wire3(105);
	sub_wire1(5, 106)    <= sub_wire3(106);
	sub_wire1(5, 107)    <= sub_wire3(107);
	sub_wire1(5, 108)    <= sub_wire3(108);
	sub_wire1(5, 109)    <= sub_wire3(109);
	sub_wire1(5, 110)    <= sub_wire3(110);
	sub_wire1(5, 111)    <= sub_wire3(111);
	sub_wire1(5, 112)    <= sub_wire3(112);
	sub_wire1(5, 113)    <= sub_wire3(113);
	sub_wire1(5, 114)    <= sub_wire3(114);
	sub_wire1(5, 115)    <= sub_wire3(115);
	sub_wire1(5, 116)    <= sub_wire3(116);
	sub_wire1(5, 117)    <= sub_wire3(117);
	sub_wire1(5, 118)    <= sub_wire3(118);
	sub_wire1(5, 119)    <= sub_wire3(119);
	sub_wire1(5, 120)    <= sub_wire3(120);
	sub_wire1(5, 121)    <= sub_wire3(121);
	sub_wire1(5, 122)    <= sub_wire3(122);
	sub_wire1(5, 123)    <= sub_wire3(123);
	sub_wire1(5, 124)    <= sub_wire3(124);
	sub_wire1(5, 125)    <= sub_wire3(125);
	sub_wire1(5, 126)    <= sub_wire3(126);
	sub_wire1(5, 127)    <= sub_wire3(127);
	sub_wire1(5, 128)    <= sub_wire3(128);
	sub_wire1(5, 129)    <= sub_wire3(129);
	sub_wire1(5, 130)    <= sub_wire3(130);
	sub_wire1(5, 131)    <= sub_wire3(131);
	sub_wire1(5, 132)    <= sub_wire3(132);
	sub_wire1(5, 133)    <= sub_wire3(133);
	sub_wire1(5, 134)    <= sub_wire3(134);
	sub_wire1(5, 135)    <= sub_wire3(135);
	sub_wire1(5, 136)    <= sub_wire3(136);
	sub_wire1(5, 137)    <= sub_wire3(137);
	sub_wire1(5, 138)    <= sub_wire3(138);
	sub_wire1(5, 139)    <= sub_wire3(139);
	sub_wire1(5, 140)    <= sub_wire3(140);
	sub_wire1(5, 141)    <= sub_wire3(141);
	sub_wire1(5, 142)    <= sub_wire3(142);
	sub_wire1(5, 143)    <= sub_wire3(143);
	sub_wire1(5, 144)    <= sub_wire3(144);
	sub_wire1(5, 145)    <= sub_wire3(145);
	sub_wire1(5, 146)    <= sub_wire3(146);
	sub_wire1(5, 147)    <= sub_wire3(147);
	sub_wire1(5, 148)    <= sub_wire3(148);
	sub_wire1(5, 149)    <= sub_wire3(149);
	sub_wire1(5, 150)    <= sub_wire3(150);
	sub_wire1(5, 151)    <= sub_wire3(151);
	sub_wire1(5, 152)    <= sub_wire3(152);
	sub_wire1(5, 153)    <= sub_wire3(153);
	sub_wire1(5, 154)    <= sub_wire3(154);
	sub_wire1(5, 155)    <= sub_wire3(155);
	sub_wire1(5, 156)    <= sub_wire3(156);
	sub_wire1(5, 157)    <= sub_wire3(157);
	sub_wire1(5, 158)    <= sub_wire3(158);
	sub_wire1(5, 159)    <= sub_wire3(159);
	sub_wire1(5, 160)    <= sub_wire3(160);
	sub_wire1(5, 161)    <= sub_wire3(161);
	sub_wire1(5, 162)    <= sub_wire3(162);
	sub_wire1(5, 163)    <= sub_wire3(163);
	sub_wire1(5, 164)    <= sub_wire3(164);
	sub_wire1(5, 165)    <= sub_wire3(165);
	sub_wire1(5, 166)    <= sub_wire3(166);
	sub_wire1(5, 167)    <= sub_wire3(167);
	sub_wire1(5, 168)    <= sub_wire3(168);
	sub_wire1(5, 169)    <= sub_wire3(169);
	sub_wire1(5, 170)    <= sub_wire3(170);
	sub_wire1(5, 171)    <= sub_wire3(171);
	sub_wire1(5, 172)    <= sub_wire3(172);
	sub_wire1(5, 173)    <= sub_wire3(173);
	sub_wire1(5, 174)    <= sub_wire3(174);
	sub_wire1(5, 175)    <= sub_wire3(175);
	sub_wire1(5, 176)    <= sub_wire3(176);
	sub_wire1(5, 177)    <= sub_wire3(177);
	sub_wire1(5, 178)    <= sub_wire3(178);
	sub_wire1(5, 179)    <= sub_wire3(179);
	sub_wire1(5, 180)    <= sub_wire3(180);
	sub_wire1(5, 181)    <= sub_wire3(181);
	sub_wire1(5, 182)    <= sub_wire3(182);
	sub_wire1(5, 183)    <= sub_wire3(183);
	sub_wire1(5, 184)    <= sub_wire3(184);
	sub_wire1(5, 185)    <= sub_wire3(185);
	sub_wire1(5, 186)    <= sub_wire3(186);
	sub_wire1(5, 187)    <= sub_wire3(187);
	sub_wire1(5, 188)    <= sub_wire3(188);
	sub_wire1(5, 189)    <= sub_wire3(189);
	sub_wire1(5, 190)    <= sub_wire3(190);
	sub_wire1(5, 191)    <= sub_wire3(191);
	sub_wire1(5, 192)    <= sub_wire3(192);
	sub_wire1(5, 193)    <= sub_wire3(193);
	sub_wire1(5, 194)    <= sub_wire3(194);
	sub_wire1(5, 195)    <= sub_wire3(195);
	sub_wire1(5, 196)    <= sub_wire3(196);
	sub_wire1(5, 197)    <= sub_wire3(197);
	sub_wire1(5, 198)    <= sub_wire3(198);
	sub_wire1(5, 199)    <= sub_wire3(199);
	sub_wire1(5, 200)    <= sub_wire3(200);
	sub_wire1(5, 201)    <= sub_wire3(201);
	sub_wire1(5, 202)    <= sub_wire3(202);
	sub_wire1(5, 203)    <= sub_wire3(203);
	sub_wire1(5, 204)    <= sub_wire3(204);
	sub_wire1(5, 205)    <= sub_wire3(205);
	sub_wire1(5, 206)    <= sub_wire3(206);
	sub_wire1(5, 207)    <= sub_wire3(207);
	sub_wire1(5, 208)    <= sub_wire3(208);
	sub_wire1(5, 209)    <= sub_wire3(209);
	sub_wire1(5, 210)    <= sub_wire3(210);
	sub_wire1(5, 211)    <= sub_wire3(211);
	sub_wire1(5, 212)    <= sub_wire3(212);
	sub_wire1(5, 213)    <= sub_wire3(213);
	sub_wire1(5, 214)    <= sub_wire3(214);
	sub_wire1(5, 215)    <= sub_wire3(215);
	sub_wire1(5, 216)    <= sub_wire3(216);
	sub_wire1(5, 217)    <= sub_wire3(217);
	sub_wire1(5, 218)    <= sub_wire3(218);
	sub_wire1(5, 219)    <= sub_wire3(219);
	sub_wire1(5, 220)    <= sub_wire3(220);
	sub_wire1(5, 221)    <= sub_wire3(221);
	sub_wire1(5, 222)    <= sub_wire3(222);
	sub_wire1(5, 223)    <= sub_wire3(223);
	sub_wire1(5, 224)    <= sub_wire3(224);
	sub_wire1(5, 225)    <= sub_wire3(225);
	sub_wire1(5, 226)    <= sub_wire3(226);
	sub_wire1(5, 227)    <= sub_wire3(227);
	sub_wire1(5, 228)    <= sub_wire3(228);
	sub_wire1(5, 229)    <= sub_wire3(229);
	sub_wire1(5, 230)    <= sub_wire3(230);
	sub_wire1(5, 231)    <= sub_wire3(231);
	sub_wire1(5, 232)    <= sub_wire3(232);
	sub_wire1(5, 233)    <= sub_wire3(233);
	sub_wire1(5, 234)    <= sub_wire3(234);
	sub_wire1(5, 235)    <= sub_wire3(235);
	sub_wire1(5, 236)    <= sub_wire3(236);
	sub_wire1(5, 237)    <= sub_wire3(237);
	sub_wire1(5, 238)    <= sub_wire3(238);
	sub_wire1(5, 239)    <= sub_wire3(239);
	sub_wire1(5, 240)    <= sub_wire3(240);
	sub_wire1(5, 241)    <= sub_wire3(241);
	sub_wire1(5, 242)    <= sub_wire3(242);
	sub_wire1(5, 243)    <= sub_wire3(243);
	sub_wire1(5, 244)    <= sub_wire3(244);
	sub_wire1(5, 245)    <= sub_wire3(245);
	sub_wire1(5, 246)    <= sub_wire3(246);
	sub_wire1(5, 247)    <= sub_wire3(247);
	sub_wire1(5, 248)    <= sub_wire3(248);
	sub_wire1(5, 249)    <= sub_wire3(249);
	sub_wire1(5, 250)    <= sub_wire3(250);
	sub_wire1(5, 251)    <= sub_wire3(251);
	sub_wire1(5, 252)    <= sub_wire3(252);
	sub_wire1(5, 253)    <= sub_wire3(253);
	sub_wire1(5, 254)    <= sub_wire3(254);
	sub_wire1(5, 255)    <= sub_wire3(255);
	sub_wire1(4, 0)    <= sub_wire4(0);
	sub_wire1(4, 1)    <= sub_wire4(1);
	sub_wire1(4, 2)    <= sub_wire4(2);
	sub_wire1(4, 3)    <= sub_wire4(3);
	sub_wire1(4, 4)    <= sub_wire4(4);
	sub_wire1(4, 5)    <= sub_wire4(5);
	sub_wire1(4, 6)    <= sub_wire4(6);
	sub_wire1(4, 7)    <= sub_wire4(7);
	sub_wire1(4, 8)    <= sub_wire4(8);
	sub_wire1(4, 9)    <= sub_wire4(9);
	sub_wire1(4, 10)    <= sub_wire4(10);
	sub_wire1(4, 11)    <= sub_wire4(11);
	sub_wire1(4, 12)    <= sub_wire4(12);
	sub_wire1(4, 13)    <= sub_wire4(13);
	sub_wire1(4, 14)    <= sub_wire4(14);
	sub_wire1(4, 15)    <= sub_wire4(15);
	sub_wire1(4, 16)    <= sub_wire4(16);
	sub_wire1(4, 17)    <= sub_wire4(17);
	sub_wire1(4, 18)    <= sub_wire4(18);
	sub_wire1(4, 19)    <= sub_wire4(19);
	sub_wire1(4, 20)    <= sub_wire4(20);
	sub_wire1(4, 21)    <= sub_wire4(21);
	sub_wire1(4, 22)    <= sub_wire4(22);
	sub_wire1(4, 23)    <= sub_wire4(23);
	sub_wire1(4, 24)    <= sub_wire4(24);
	sub_wire1(4, 25)    <= sub_wire4(25);
	sub_wire1(4, 26)    <= sub_wire4(26);
	sub_wire1(4, 27)    <= sub_wire4(27);
	sub_wire1(4, 28)    <= sub_wire4(28);
	sub_wire1(4, 29)    <= sub_wire4(29);
	sub_wire1(4, 30)    <= sub_wire4(30);
	sub_wire1(4, 31)    <= sub_wire4(31);
	sub_wire1(4, 32)    <= sub_wire4(32);
	sub_wire1(4, 33)    <= sub_wire4(33);
	sub_wire1(4, 34)    <= sub_wire4(34);
	sub_wire1(4, 35)    <= sub_wire4(35);
	sub_wire1(4, 36)    <= sub_wire4(36);
	sub_wire1(4, 37)    <= sub_wire4(37);
	sub_wire1(4, 38)    <= sub_wire4(38);
	sub_wire1(4, 39)    <= sub_wire4(39);
	sub_wire1(4, 40)    <= sub_wire4(40);
	sub_wire1(4, 41)    <= sub_wire4(41);
	sub_wire1(4, 42)    <= sub_wire4(42);
	sub_wire1(4, 43)    <= sub_wire4(43);
	sub_wire1(4, 44)    <= sub_wire4(44);
	sub_wire1(4, 45)    <= sub_wire4(45);
	sub_wire1(4, 46)    <= sub_wire4(46);
	sub_wire1(4, 47)    <= sub_wire4(47);
	sub_wire1(4, 48)    <= sub_wire4(48);
	sub_wire1(4, 49)    <= sub_wire4(49);
	sub_wire1(4, 50)    <= sub_wire4(50);
	sub_wire1(4, 51)    <= sub_wire4(51);
	sub_wire1(4, 52)    <= sub_wire4(52);
	sub_wire1(4, 53)    <= sub_wire4(53);
	sub_wire1(4, 54)    <= sub_wire4(54);
	sub_wire1(4, 55)    <= sub_wire4(55);
	sub_wire1(4, 56)    <= sub_wire4(56);
	sub_wire1(4, 57)    <= sub_wire4(57);
	sub_wire1(4, 58)    <= sub_wire4(58);
	sub_wire1(4, 59)    <= sub_wire4(59);
	sub_wire1(4, 60)    <= sub_wire4(60);
	sub_wire1(4, 61)    <= sub_wire4(61);
	sub_wire1(4, 62)    <= sub_wire4(62);
	sub_wire1(4, 63)    <= sub_wire4(63);
	sub_wire1(4, 64)    <= sub_wire4(64);
	sub_wire1(4, 65)    <= sub_wire4(65);
	sub_wire1(4, 66)    <= sub_wire4(66);
	sub_wire1(4, 67)    <= sub_wire4(67);
	sub_wire1(4, 68)    <= sub_wire4(68);
	sub_wire1(4, 69)    <= sub_wire4(69);
	sub_wire1(4, 70)    <= sub_wire4(70);
	sub_wire1(4, 71)    <= sub_wire4(71);
	sub_wire1(4, 72)    <= sub_wire4(72);
	sub_wire1(4, 73)    <= sub_wire4(73);
	sub_wire1(4, 74)    <= sub_wire4(74);
	sub_wire1(4, 75)    <= sub_wire4(75);
	sub_wire1(4, 76)    <= sub_wire4(76);
	sub_wire1(4, 77)    <= sub_wire4(77);
	sub_wire1(4, 78)    <= sub_wire4(78);
	sub_wire1(4, 79)    <= sub_wire4(79);
	sub_wire1(4, 80)    <= sub_wire4(80);
	sub_wire1(4, 81)    <= sub_wire4(81);
	sub_wire1(4, 82)    <= sub_wire4(82);
	sub_wire1(4, 83)    <= sub_wire4(83);
	sub_wire1(4, 84)    <= sub_wire4(84);
	sub_wire1(4, 85)    <= sub_wire4(85);
	sub_wire1(4, 86)    <= sub_wire4(86);
	sub_wire1(4, 87)    <= sub_wire4(87);
	sub_wire1(4, 88)    <= sub_wire4(88);
	sub_wire1(4, 89)    <= sub_wire4(89);
	sub_wire1(4, 90)    <= sub_wire4(90);
	sub_wire1(4, 91)    <= sub_wire4(91);
	sub_wire1(4, 92)    <= sub_wire4(92);
	sub_wire1(4, 93)    <= sub_wire4(93);
	sub_wire1(4, 94)    <= sub_wire4(94);
	sub_wire1(4, 95)    <= sub_wire4(95);
	sub_wire1(4, 96)    <= sub_wire4(96);
	sub_wire1(4, 97)    <= sub_wire4(97);
	sub_wire1(4, 98)    <= sub_wire4(98);
	sub_wire1(4, 99)    <= sub_wire4(99);
	sub_wire1(4, 100)    <= sub_wire4(100);
	sub_wire1(4, 101)    <= sub_wire4(101);
	sub_wire1(4, 102)    <= sub_wire4(102);
	sub_wire1(4, 103)    <= sub_wire4(103);
	sub_wire1(4, 104)    <= sub_wire4(104);
	sub_wire1(4, 105)    <= sub_wire4(105);
	sub_wire1(4, 106)    <= sub_wire4(106);
	sub_wire1(4, 107)    <= sub_wire4(107);
	sub_wire1(4, 108)    <= sub_wire4(108);
	sub_wire1(4, 109)    <= sub_wire4(109);
	sub_wire1(4, 110)    <= sub_wire4(110);
	sub_wire1(4, 111)    <= sub_wire4(111);
	sub_wire1(4, 112)    <= sub_wire4(112);
	sub_wire1(4, 113)    <= sub_wire4(113);
	sub_wire1(4, 114)    <= sub_wire4(114);
	sub_wire1(4, 115)    <= sub_wire4(115);
	sub_wire1(4, 116)    <= sub_wire4(116);
	sub_wire1(4, 117)    <= sub_wire4(117);
	sub_wire1(4, 118)    <= sub_wire4(118);
	sub_wire1(4, 119)    <= sub_wire4(119);
	sub_wire1(4, 120)    <= sub_wire4(120);
	sub_wire1(4, 121)    <= sub_wire4(121);
	sub_wire1(4, 122)    <= sub_wire4(122);
	sub_wire1(4, 123)    <= sub_wire4(123);
	sub_wire1(4, 124)    <= sub_wire4(124);
	sub_wire1(4, 125)    <= sub_wire4(125);
	sub_wire1(4, 126)    <= sub_wire4(126);
	sub_wire1(4, 127)    <= sub_wire4(127);
	sub_wire1(4, 128)    <= sub_wire4(128);
	sub_wire1(4, 129)    <= sub_wire4(129);
	sub_wire1(4, 130)    <= sub_wire4(130);
	sub_wire1(4, 131)    <= sub_wire4(131);
	sub_wire1(4, 132)    <= sub_wire4(132);
	sub_wire1(4, 133)    <= sub_wire4(133);
	sub_wire1(4, 134)    <= sub_wire4(134);
	sub_wire1(4, 135)    <= sub_wire4(135);
	sub_wire1(4, 136)    <= sub_wire4(136);
	sub_wire1(4, 137)    <= sub_wire4(137);
	sub_wire1(4, 138)    <= sub_wire4(138);
	sub_wire1(4, 139)    <= sub_wire4(139);
	sub_wire1(4, 140)    <= sub_wire4(140);
	sub_wire1(4, 141)    <= sub_wire4(141);
	sub_wire1(4, 142)    <= sub_wire4(142);
	sub_wire1(4, 143)    <= sub_wire4(143);
	sub_wire1(4, 144)    <= sub_wire4(144);
	sub_wire1(4, 145)    <= sub_wire4(145);
	sub_wire1(4, 146)    <= sub_wire4(146);
	sub_wire1(4, 147)    <= sub_wire4(147);
	sub_wire1(4, 148)    <= sub_wire4(148);
	sub_wire1(4, 149)    <= sub_wire4(149);
	sub_wire1(4, 150)    <= sub_wire4(150);
	sub_wire1(4, 151)    <= sub_wire4(151);
	sub_wire1(4, 152)    <= sub_wire4(152);
	sub_wire1(4, 153)    <= sub_wire4(153);
	sub_wire1(4, 154)    <= sub_wire4(154);
	sub_wire1(4, 155)    <= sub_wire4(155);
	sub_wire1(4, 156)    <= sub_wire4(156);
	sub_wire1(4, 157)    <= sub_wire4(157);
	sub_wire1(4, 158)    <= sub_wire4(158);
	sub_wire1(4, 159)    <= sub_wire4(159);
	sub_wire1(4, 160)    <= sub_wire4(160);
	sub_wire1(4, 161)    <= sub_wire4(161);
	sub_wire1(4, 162)    <= sub_wire4(162);
	sub_wire1(4, 163)    <= sub_wire4(163);
	sub_wire1(4, 164)    <= sub_wire4(164);
	sub_wire1(4, 165)    <= sub_wire4(165);
	sub_wire1(4, 166)    <= sub_wire4(166);
	sub_wire1(4, 167)    <= sub_wire4(167);
	sub_wire1(4, 168)    <= sub_wire4(168);
	sub_wire1(4, 169)    <= sub_wire4(169);
	sub_wire1(4, 170)    <= sub_wire4(170);
	sub_wire1(4, 171)    <= sub_wire4(171);
	sub_wire1(4, 172)    <= sub_wire4(172);
	sub_wire1(4, 173)    <= sub_wire4(173);
	sub_wire1(4, 174)    <= sub_wire4(174);
	sub_wire1(4, 175)    <= sub_wire4(175);
	sub_wire1(4, 176)    <= sub_wire4(176);
	sub_wire1(4, 177)    <= sub_wire4(177);
	sub_wire1(4, 178)    <= sub_wire4(178);
	sub_wire1(4, 179)    <= sub_wire4(179);
	sub_wire1(4, 180)    <= sub_wire4(180);
	sub_wire1(4, 181)    <= sub_wire4(181);
	sub_wire1(4, 182)    <= sub_wire4(182);
	sub_wire1(4, 183)    <= sub_wire4(183);
	sub_wire1(4, 184)    <= sub_wire4(184);
	sub_wire1(4, 185)    <= sub_wire4(185);
	sub_wire1(4, 186)    <= sub_wire4(186);
	sub_wire1(4, 187)    <= sub_wire4(187);
	sub_wire1(4, 188)    <= sub_wire4(188);
	sub_wire1(4, 189)    <= sub_wire4(189);
	sub_wire1(4, 190)    <= sub_wire4(190);
	sub_wire1(4, 191)    <= sub_wire4(191);
	sub_wire1(4, 192)    <= sub_wire4(192);
	sub_wire1(4, 193)    <= sub_wire4(193);
	sub_wire1(4, 194)    <= sub_wire4(194);
	sub_wire1(4, 195)    <= sub_wire4(195);
	sub_wire1(4, 196)    <= sub_wire4(196);
	sub_wire1(4, 197)    <= sub_wire4(197);
	sub_wire1(4, 198)    <= sub_wire4(198);
	sub_wire1(4, 199)    <= sub_wire4(199);
	sub_wire1(4, 200)    <= sub_wire4(200);
	sub_wire1(4, 201)    <= sub_wire4(201);
	sub_wire1(4, 202)    <= sub_wire4(202);
	sub_wire1(4, 203)    <= sub_wire4(203);
	sub_wire1(4, 204)    <= sub_wire4(204);
	sub_wire1(4, 205)    <= sub_wire4(205);
	sub_wire1(4, 206)    <= sub_wire4(206);
	sub_wire1(4, 207)    <= sub_wire4(207);
	sub_wire1(4, 208)    <= sub_wire4(208);
	sub_wire1(4, 209)    <= sub_wire4(209);
	sub_wire1(4, 210)    <= sub_wire4(210);
	sub_wire1(4, 211)    <= sub_wire4(211);
	sub_wire1(4, 212)    <= sub_wire4(212);
	sub_wire1(4, 213)    <= sub_wire4(213);
	sub_wire1(4, 214)    <= sub_wire4(214);
	sub_wire1(4, 215)    <= sub_wire4(215);
	sub_wire1(4, 216)    <= sub_wire4(216);
	sub_wire1(4, 217)    <= sub_wire4(217);
	sub_wire1(4, 218)    <= sub_wire4(218);
	sub_wire1(4, 219)    <= sub_wire4(219);
	sub_wire1(4, 220)    <= sub_wire4(220);
	sub_wire1(4, 221)    <= sub_wire4(221);
	sub_wire1(4, 222)    <= sub_wire4(222);
	sub_wire1(4, 223)    <= sub_wire4(223);
	sub_wire1(4, 224)    <= sub_wire4(224);
	sub_wire1(4, 225)    <= sub_wire4(225);
	sub_wire1(4, 226)    <= sub_wire4(226);
	sub_wire1(4, 227)    <= sub_wire4(227);
	sub_wire1(4, 228)    <= sub_wire4(228);
	sub_wire1(4, 229)    <= sub_wire4(229);
	sub_wire1(4, 230)    <= sub_wire4(230);
	sub_wire1(4, 231)    <= sub_wire4(231);
	sub_wire1(4, 232)    <= sub_wire4(232);
	sub_wire1(4, 233)    <= sub_wire4(233);
	sub_wire1(4, 234)    <= sub_wire4(234);
	sub_wire1(4, 235)    <= sub_wire4(235);
	sub_wire1(4, 236)    <= sub_wire4(236);
	sub_wire1(4, 237)    <= sub_wire4(237);
	sub_wire1(4, 238)    <= sub_wire4(238);
	sub_wire1(4, 239)    <= sub_wire4(239);
	sub_wire1(4, 240)    <= sub_wire4(240);
	sub_wire1(4, 241)    <= sub_wire4(241);
	sub_wire1(4, 242)    <= sub_wire4(242);
	sub_wire1(4, 243)    <= sub_wire4(243);
	sub_wire1(4, 244)    <= sub_wire4(244);
	sub_wire1(4, 245)    <= sub_wire4(245);
	sub_wire1(4, 246)    <= sub_wire4(246);
	sub_wire1(4, 247)    <= sub_wire4(247);
	sub_wire1(4, 248)    <= sub_wire4(248);
	sub_wire1(4, 249)    <= sub_wire4(249);
	sub_wire1(4, 250)    <= sub_wire4(250);
	sub_wire1(4, 251)    <= sub_wire4(251);
	sub_wire1(4, 252)    <= sub_wire4(252);
	sub_wire1(4, 253)    <= sub_wire4(253);
	sub_wire1(4, 254)    <= sub_wire4(254);
	sub_wire1(4, 255)    <= sub_wire4(255);
	sub_wire1(3, 0)    <= sub_wire5(0);
	sub_wire1(3, 1)    <= sub_wire5(1);
	sub_wire1(3, 2)    <= sub_wire5(2);
	sub_wire1(3, 3)    <= sub_wire5(3);
	sub_wire1(3, 4)    <= sub_wire5(4);
	sub_wire1(3, 5)    <= sub_wire5(5);
	sub_wire1(3, 6)    <= sub_wire5(6);
	sub_wire1(3, 7)    <= sub_wire5(7);
	sub_wire1(3, 8)    <= sub_wire5(8);
	sub_wire1(3, 9)    <= sub_wire5(9);
	sub_wire1(3, 10)    <= sub_wire5(10);
	sub_wire1(3, 11)    <= sub_wire5(11);
	sub_wire1(3, 12)    <= sub_wire5(12);
	sub_wire1(3, 13)    <= sub_wire5(13);
	sub_wire1(3, 14)    <= sub_wire5(14);
	sub_wire1(3, 15)    <= sub_wire5(15);
	sub_wire1(3, 16)    <= sub_wire5(16);
	sub_wire1(3, 17)    <= sub_wire5(17);
	sub_wire1(3, 18)    <= sub_wire5(18);
	sub_wire1(3, 19)    <= sub_wire5(19);
	sub_wire1(3, 20)    <= sub_wire5(20);
	sub_wire1(3, 21)    <= sub_wire5(21);
	sub_wire1(3, 22)    <= sub_wire5(22);
	sub_wire1(3, 23)    <= sub_wire5(23);
	sub_wire1(3, 24)    <= sub_wire5(24);
	sub_wire1(3, 25)    <= sub_wire5(25);
	sub_wire1(3, 26)    <= sub_wire5(26);
	sub_wire1(3, 27)    <= sub_wire5(27);
	sub_wire1(3, 28)    <= sub_wire5(28);
	sub_wire1(3, 29)    <= sub_wire5(29);
	sub_wire1(3, 30)    <= sub_wire5(30);
	sub_wire1(3, 31)    <= sub_wire5(31);
	sub_wire1(3, 32)    <= sub_wire5(32);
	sub_wire1(3, 33)    <= sub_wire5(33);
	sub_wire1(3, 34)    <= sub_wire5(34);
	sub_wire1(3, 35)    <= sub_wire5(35);
	sub_wire1(3, 36)    <= sub_wire5(36);
	sub_wire1(3, 37)    <= sub_wire5(37);
	sub_wire1(3, 38)    <= sub_wire5(38);
	sub_wire1(3, 39)    <= sub_wire5(39);
	sub_wire1(3, 40)    <= sub_wire5(40);
	sub_wire1(3, 41)    <= sub_wire5(41);
	sub_wire1(3, 42)    <= sub_wire5(42);
	sub_wire1(3, 43)    <= sub_wire5(43);
	sub_wire1(3, 44)    <= sub_wire5(44);
	sub_wire1(3, 45)    <= sub_wire5(45);
	sub_wire1(3, 46)    <= sub_wire5(46);
	sub_wire1(3, 47)    <= sub_wire5(47);
	sub_wire1(3, 48)    <= sub_wire5(48);
	sub_wire1(3, 49)    <= sub_wire5(49);
	sub_wire1(3, 50)    <= sub_wire5(50);
	sub_wire1(3, 51)    <= sub_wire5(51);
	sub_wire1(3, 52)    <= sub_wire5(52);
	sub_wire1(3, 53)    <= sub_wire5(53);
	sub_wire1(3, 54)    <= sub_wire5(54);
	sub_wire1(3, 55)    <= sub_wire5(55);
	sub_wire1(3, 56)    <= sub_wire5(56);
	sub_wire1(3, 57)    <= sub_wire5(57);
	sub_wire1(3, 58)    <= sub_wire5(58);
	sub_wire1(3, 59)    <= sub_wire5(59);
	sub_wire1(3, 60)    <= sub_wire5(60);
	sub_wire1(3, 61)    <= sub_wire5(61);
	sub_wire1(3, 62)    <= sub_wire5(62);
	sub_wire1(3, 63)    <= sub_wire5(63);
	sub_wire1(3, 64)    <= sub_wire5(64);
	sub_wire1(3, 65)    <= sub_wire5(65);
	sub_wire1(3, 66)    <= sub_wire5(66);
	sub_wire1(3, 67)    <= sub_wire5(67);
	sub_wire1(3, 68)    <= sub_wire5(68);
	sub_wire1(3, 69)    <= sub_wire5(69);
	sub_wire1(3, 70)    <= sub_wire5(70);
	sub_wire1(3, 71)    <= sub_wire5(71);
	sub_wire1(3, 72)    <= sub_wire5(72);
	sub_wire1(3, 73)    <= sub_wire5(73);
	sub_wire1(3, 74)    <= sub_wire5(74);
	sub_wire1(3, 75)    <= sub_wire5(75);
	sub_wire1(3, 76)    <= sub_wire5(76);
	sub_wire1(3, 77)    <= sub_wire5(77);
	sub_wire1(3, 78)    <= sub_wire5(78);
	sub_wire1(3, 79)    <= sub_wire5(79);
	sub_wire1(3, 80)    <= sub_wire5(80);
	sub_wire1(3, 81)    <= sub_wire5(81);
	sub_wire1(3, 82)    <= sub_wire5(82);
	sub_wire1(3, 83)    <= sub_wire5(83);
	sub_wire1(3, 84)    <= sub_wire5(84);
	sub_wire1(3, 85)    <= sub_wire5(85);
	sub_wire1(3, 86)    <= sub_wire5(86);
	sub_wire1(3, 87)    <= sub_wire5(87);
	sub_wire1(3, 88)    <= sub_wire5(88);
	sub_wire1(3, 89)    <= sub_wire5(89);
	sub_wire1(3, 90)    <= sub_wire5(90);
	sub_wire1(3, 91)    <= sub_wire5(91);
	sub_wire1(3, 92)    <= sub_wire5(92);
	sub_wire1(3, 93)    <= sub_wire5(93);
	sub_wire1(3, 94)    <= sub_wire5(94);
	sub_wire1(3, 95)    <= sub_wire5(95);
	sub_wire1(3, 96)    <= sub_wire5(96);
	sub_wire1(3, 97)    <= sub_wire5(97);
	sub_wire1(3, 98)    <= sub_wire5(98);
	sub_wire1(3, 99)    <= sub_wire5(99);
	sub_wire1(3, 100)    <= sub_wire5(100);
	sub_wire1(3, 101)    <= sub_wire5(101);
	sub_wire1(3, 102)    <= sub_wire5(102);
	sub_wire1(3, 103)    <= sub_wire5(103);
	sub_wire1(3, 104)    <= sub_wire5(104);
	sub_wire1(3, 105)    <= sub_wire5(105);
	sub_wire1(3, 106)    <= sub_wire5(106);
	sub_wire1(3, 107)    <= sub_wire5(107);
	sub_wire1(3, 108)    <= sub_wire5(108);
	sub_wire1(3, 109)    <= sub_wire5(109);
	sub_wire1(3, 110)    <= sub_wire5(110);
	sub_wire1(3, 111)    <= sub_wire5(111);
	sub_wire1(3, 112)    <= sub_wire5(112);
	sub_wire1(3, 113)    <= sub_wire5(113);
	sub_wire1(3, 114)    <= sub_wire5(114);
	sub_wire1(3, 115)    <= sub_wire5(115);
	sub_wire1(3, 116)    <= sub_wire5(116);
	sub_wire1(3, 117)    <= sub_wire5(117);
	sub_wire1(3, 118)    <= sub_wire5(118);
	sub_wire1(3, 119)    <= sub_wire5(119);
	sub_wire1(3, 120)    <= sub_wire5(120);
	sub_wire1(3, 121)    <= sub_wire5(121);
	sub_wire1(3, 122)    <= sub_wire5(122);
	sub_wire1(3, 123)    <= sub_wire5(123);
	sub_wire1(3, 124)    <= sub_wire5(124);
	sub_wire1(3, 125)    <= sub_wire5(125);
	sub_wire1(3, 126)    <= sub_wire5(126);
	sub_wire1(3, 127)    <= sub_wire5(127);
	sub_wire1(3, 128)    <= sub_wire5(128);
	sub_wire1(3, 129)    <= sub_wire5(129);
	sub_wire1(3, 130)    <= sub_wire5(130);
	sub_wire1(3, 131)    <= sub_wire5(131);
	sub_wire1(3, 132)    <= sub_wire5(132);
	sub_wire1(3, 133)    <= sub_wire5(133);
	sub_wire1(3, 134)    <= sub_wire5(134);
	sub_wire1(3, 135)    <= sub_wire5(135);
	sub_wire1(3, 136)    <= sub_wire5(136);
	sub_wire1(3, 137)    <= sub_wire5(137);
	sub_wire1(3, 138)    <= sub_wire5(138);
	sub_wire1(3, 139)    <= sub_wire5(139);
	sub_wire1(3, 140)    <= sub_wire5(140);
	sub_wire1(3, 141)    <= sub_wire5(141);
	sub_wire1(3, 142)    <= sub_wire5(142);
	sub_wire1(3, 143)    <= sub_wire5(143);
	sub_wire1(3, 144)    <= sub_wire5(144);
	sub_wire1(3, 145)    <= sub_wire5(145);
	sub_wire1(3, 146)    <= sub_wire5(146);
	sub_wire1(3, 147)    <= sub_wire5(147);
	sub_wire1(3, 148)    <= sub_wire5(148);
	sub_wire1(3, 149)    <= sub_wire5(149);
	sub_wire1(3, 150)    <= sub_wire5(150);
	sub_wire1(3, 151)    <= sub_wire5(151);
	sub_wire1(3, 152)    <= sub_wire5(152);
	sub_wire1(3, 153)    <= sub_wire5(153);
	sub_wire1(3, 154)    <= sub_wire5(154);
	sub_wire1(3, 155)    <= sub_wire5(155);
	sub_wire1(3, 156)    <= sub_wire5(156);
	sub_wire1(3, 157)    <= sub_wire5(157);
	sub_wire1(3, 158)    <= sub_wire5(158);
	sub_wire1(3, 159)    <= sub_wire5(159);
	sub_wire1(3, 160)    <= sub_wire5(160);
	sub_wire1(3, 161)    <= sub_wire5(161);
	sub_wire1(3, 162)    <= sub_wire5(162);
	sub_wire1(3, 163)    <= sub_wire5(163);
	sub_wire1(3, 164)    <= sub_wire5(164);
	sub_wire1(3, 165)    <= sub_wire5(165);
	sub_wire1(3, 166)    <= sub_wire5(166);
	sub_wire1(3, 167)    <= sub_wire5(167);
	sub_wire1(3, 168)    <= sub_wire5(168);
	sub_wire1(3, 169)    <= sub_wire5(169);
	sub_wire1(3, 170)    <= sub_wire5(170);
	sub_wire1(3, 171)    <= sub_wire5(171);
	sub_wire1(3, 172)    <= sub_wire5(172);
	sub_wire1(3, 173)    <= sub_wire5(173);
	sub_wire1(3, 174)    <= sub_wire5(174);
	sub_wire1(3, 175)    <= sub_wire5(175);
	sub_wire1(3, 176)    <= sub_wire5(176);
	sub_wire1(3, 177)    <= sub_wire5(177);
	sub_wire1(3, 178)    <= sub_wire5(178);
	sub_wire1(3, 179)    <= sub_wire5(179);
	sub_wire1(3, 180)    <= sub_wire5(180);
	sub_wire1(3, 181)    <= sub_wire5(181);
	sub_wire1(3, 182)    <= sub_wire5(182);
	sub_wire1(3, 183)    <= sub_wire5(183);
	sub_wire1(3, 184)    <= sub_wire5(184);
	sub_wire1(3, 185)    <= sub_wire5(185);
	sub_wire1(3, 186)    <= sub_wire5(186);
	sub_wire1(3, 187)    <= sub_wire5(187);
	sub_wire1(3, 188)    <= sub_wire5(188);
	sub_wire1(3, 189)    <= sub_wire5(189);
	sub_wire1(3, 190)    <= sub_wire5(190);
	sub_wire1(3, 191)    <= sub_wire5(191);
	sub_wire1(3, 192)    <= sub_wire5(192);
	sub_wire1(3, 193)    <= sub_wire5(193);
	sub_wire1(3, 194)    <= sub_wire5(194);
	sub_wire1(3, 195)    <= sub_wire5(195);
	sub_wire1(3, 196)    <= sub_wire5(196);
	sub_wire1(3, 197)    <= sub_wire5(197);
	sub_wire1(3, 198)    <= sub_wire5(198);
	sub_wire1(3, 199)    <= sub_wire5(199);
	sub_wire1(3, 200)    <= sub_wire5(200);
	sub_wire1(3, 201)    <= sub_wire5(201);
	sub_wire1(3, 202)    <= sub_wire5(202);
	sub_wire1(3, 203)    <= sub_wire5(203);
	sub_wire1(3, 204)    <= sub_wire5(204);
	sub_wire1(3, 205)    <= sub_wire5(205);
	sub_wire1(3, 206)    <= sub_wire5(206);
	sub_wire1(3, 207)    <= sub_wire5(207);
	sub_wire1(3, 208)    <= sub_wire5(208);
	sub_wire1(3, 209)    <= sub_wire5(209);
	sub_wire1(3, 210)    <= sub_wire5(210);
	sub_wire1(3, 211)    <= sub_wire5(211);
	sub_wire1(3, 212)    <= sub_wire5(212);
	sub_wire1(3, 213)    <= sub_wire5(213);
	sub_wire1(3, 214)    <= sub_wire5(214);
	sub_wire1(3, 215)    <= sub_wire5(215);
	sub_wire1(3, 216)    <= sub_wire5(216);
	sub_wire1(3, 217)    <= sub_wire5(217);
	sub_wire1(3, 218)    <= sub_wire5(218);
	sub_wire1(3, 219)    <= sub_wire5(219);
	sub_wire1(3, 220)    <= sub_wire5(220);
	sub_wire1(3, 221)    <= sub_wire5(221);
	sub_wire1(3, 222)    <= sub_wire5(222);
	sub_wire1(3, 223)    <= sub_wire5(223);
	sub_wire1(3, 224)    <= sub_wire5(224);
	sub_wire1(3, 225)    <= sub_wire5(225);
	sub_wire1(3, 226)    <= sub_wire5(226);
	sub_wire1(3, 227)    <= sub_wire5(227);
	sub_wire1(3, 228)    <= sub_wire5(228);
	sub_wire1(3, 229)    <= sub_wire5(229);
	sub_wire1(3, 230)    <= sub_wire5(230);
	sub_wire1(3, 231)    <= sub_wire5(231);
	sub_wire1(3, 232)    <= sub_wire5(232);
	sub_wire1(3, 233)    <= sub_wire5(233);
	sub_wire1(3, 234)    <= sub_wire5(234);
	sub_wire1(3, 235)    <= sub_wire5(235);
	sub_wire1(3, 236)    <= sub_wire5(236);
	sub_wire1(3, 237)    <= sub_wire5(237);
	sub_wire1(3, 238)    <= sub_wire5(238);
	sub_wire1(3, 239)    <= sub_wire5(239);
	sub_wire1(3, 240)    <= sub_wire5(240);
	sub_wire1(3, 241)    <= sub_wire5(241);
	sub_wire1(3, 242)    <= sub_wire5(242);
	sub_wire1(3, 243)    <= sub_wire5(243);
	sub_wire1(3, 244)    <= sub_wire5(244);
	sub_wire1(3, 245)    <= sub_wire5(245);
	sub_wire1(3, 246)    <= sub_wire5(246);
	sub_wire1(3, 247)    <= sub_wire5(247);
	sub_wire1(3, 248)    <= sub_wire5(248);
	sub_wire1(3, 249)    <= sub_wire5(249);
	sub_wire1(3, 250)    <= sub_wire5(250);
	sub_wire1(3, 251)    <= sub_wire5(251);
	sub_wire1(3, 252)    <= sub_wire5(252);
	sub_wire1(3, 253)    <= sub_wire5(253);
	sub_wire1(3, 254)    <= sub_wire5(254);
	sub_wire1(3, 255)    <= sub_wire5(255);
	sub_wire1(2, 0)    <= sub_wire6(0);
	sub_wire1(2, 1)    <= sub_wire6(1);
	sub_wire1(2, 2)    <= sub_wire6(2);
	sub_wire1(2, 3)    <= sub_wire6(3);
	sub_wire1(2, 4)    <= sub_wire6(4);
	sub_wire1(2, 5)    <= sub_wire6(5);
	sub_wire1(2, 6)    <= sub_wire6(6);
	sub_wire1(2, 7)    <= sub_wire6(7);
	sub_wire1(2, 8)    <= sub_wire6(8);
	sub_wire1(2, 9)    <= sub_wire6(9);
	sub_wire1(2, 10)    <= sub_wire6(10);
	sub_wire1(2, 11)    <= sub_wire6(11);
	sub_wire1(2, 12)    <= sub_wire6(12);
	sub_wire1(2, 13)    <= sub_wire6(13);
	sub_wire1(2, 14)    <= sub_wire6(14);
	sub_wire1(2, 15)    <= sub_wire6(15);
	sub_wire1(2, 16)    <= sub_wire6(16);
	sub_wire1(2, 17)    <= sub_wire6(17);
	sub_wire1(2, 18)    <= sub_wire6(18);
	sub_wire1(2, 19)    <= sub_wire6(19);
	sub_wire1(2, 20)    <= sub_wire6(20);
	sub_wire1(2, 21)    <= sub_wire6(21);
	sub_wire1(2, 22)    <= sub_wire6(22);
	sub_wire1(2, 23)    <= sub_wire6(23);
	sub_wire1(2, 24)    <= sub_wire6(24);
	sub_wire1(2, 25)    <= sub_wire6(25);
	sub_wire1(2, 26)    <= sub_wire6(26);
	sub_wire1(2, 27)    <= sub_wire6(27);
	sub_wire1(2, 28)    <= sub_wire6(28);
	sub_wire1(2, 29)    <= sub_wire6(29);
	sub_wire1(2, 30)    <= sub_wire6(30);
	sub_wire1(2, 31)    <= sub_wire6(31);
	sub_wire1(2, 32)    <= sub_wire6(32);
	sub_wire1(2, 33)    <= sub_wire6(33);
	sub_wire1(2, 34)    <= sub_wire6(34);
	sub_wire1(2, 35)    <= sub_wire6(35);
	sub_wire1(2, 36)    <= sub_wire6(36);
	sub_wire1(2, 37)    <= sub_wire6(37);
	sub_wire1(2, 38)    <= sub_wire6(38);
	sub_wire1(2, 39)    <= sub_wire6(39);
	sub_wire1(2, 40)    <= sub_wire6(40);
	sub_wire1(2, 41)    <= sub_wire6(41);
	sub_wire1(2, 42)    <= sub_wire6(42);
	sub_wire1(2, 43)    <= sub_wire6(43);
	sub_wire1(2, 44)    <= sub_wire6(44);
	sub_wire1(2, 45)    <= sub_wire6(45);
	sub_wire1(2, 46)    <= sub_wire6(46);
	sub_wire1(2, 47)    <= sub_wire6(47);
	sub_wire1(2, 48)    <= sub_wire6(48);
	sub_wire1(2, 49)    <= sub_wire6(49);
	sub_wire1(2, 50)    <= sub_wire6(50);
	sub_wire1(2, 51)    <= sub_wire6(51);
	sub_wire1(2, 52)    <= sub_wire6(52);
	sub_wire1(2, 53)    <= sub_wire6(53);
	sub_wire1(2, 54)    <= sub_wire6(54);
	sub_wire1(2, 55)    <= sub_wire6(55);
	sub_wire1(2, 56)    <= sub_wire6(56);
	sub_wire1(2, 57)    <= sub_wire6(57);
	sub_wire1(2, 58)    <= sub_wire6(58);
	sub_wire1(2, 59)    <= sub_wire6(59);
	sub_wire1(2, 60)    <= sub_wire6(60);
	sub_wire1(2, 61)    <= sub_wire6(61);
	sub_wire1(2, 62)    <= sub_wire6(62);
	sub_wire1(2, 63)    <= sub_wire6(63);
	sub_wire1(2, 64)    <= sub_wire6(64);
	sub_wire1(2, 65)    <= sub_wire6(65);
	sub_wire1(2, 66)    <= sub_wire6(66);
	sub_wire1(2, 67)    <= sub_wire6(67);
	sub_wire1(2, 68)    <= sub_wire6(68);
	sub_wire1(2, 69)    <= sub_wire6(69);
	sub_wire1(2, 70)    <= sub_wire6(70);
	sub_wire1(2, 71)    <= sub_wire6(71);
	sub_wire1(2, 72)    <= sub_wire6(72);
	sub_wire1(2, 73)    <= sub_wire6(73);
	sub_wire1(2, 74)    <= sub_wire6(74);
	sub_wire1(2, 75)    <= sub_wire6(75);
	sub_wire1(2, 76)    <= sub_wire6(76);
	sub_wire1(2, 77)    <= sub_wire6(77);
	sub_wire1(2, 78)    <= sub_wire6(78);
	sub_wire1(2, 79)    <= sub_wire6(79);
	sub_wire1(2, 80)    <= sub_wire6(80);
	sub_wire1(2, 81)    <= sub_wire6(81);
	sub_wire1(2, 82)    <= sub_wire6(82);
	sub_wire1(2, 83)    <= sub_wire6(83);
	sub_wire1(2, 84)    <= sub_wire6(84);
	sub_wire1(2, 85)    <= sub_wire6(85);
	sub_wire1(2, 86)    <= sub_wire6(86);
	sub_wire1(2, 87)    <= sub_wire6(87);
	sub_wire1(2, 88)    <= sub_wire6(88);
	sub_wire1(2, 89)    <= sub_wire6(89);
	sub_wire1(2, 90)    <= sub_wire6(90);
	sub_wire1(2, 91)    <= sub_wire6(91);
	sub_wire1(2, 92)    <= sub_wire6(92);
	sub_wire1(2, 93)    <= sub_wire6(93);
	sub_wire1(2, 94)    <= sub_wire6(94);
	sub_wire1(2, 95)    <= sub_wire6(95);
	sub_wire1(2, 96)    <= sub_wire6(96);
	sub_wire1(2, 97)    <= sub_wire6(97);
	sub_wire1(2, 98)    <= sub_wire6(98);
	sub_wire1(2, 99)    <= sub_wire6(99);
	sub_wire1(2, 100)    <= sub_wire6(100);
	sub_wire1(2, 101)    <= sub_wire6(101);
	sub_wire1(2, 102)    <= sub_wire6(102);
	sub_wire1(2, 103)    <= sub_wire6(103);
	sub_wire1(2, 104)    <= sub_wire6(104);
	sub_wire1(2, 105)    <= sub_wire6(105);
	sub_wire1(2, 106)    <= sub_wire6(106);
	sub_wire1(2, 107)    <= sub_wire6(107);
	sub_wire1(2, 108)    <= sub_wire6(108);
	sub_wire1(2, 109)    <= sub_wire6(109);
	sub_wire1(2, 110)    <= sub_wire6(110);
	sub_wire1(2, 111)    <= sub_wire6(111);
	sub_wire1(2, 112)    <= sub_wire6(112);
	sub_wire1(2, 113)    <= sub_wire6(113);
	sub_wire1(2, 114)    <= sub_wire6(114);
	sub_wire1(2, 115)    <= sub_wire6(115);
	sub_wire1(2, 116)    <= sub_wire6(116);
	sub_wire1(2, 117)    <= sub_wire6(117);
	sub_wire1(2, 118)    <= sub_wire6(118);
	sub_wire1(2, 119)    <= sub_wire6(119);
	sub_wire1(2, 120)    <= sub_wire6(120);
	sub_wire1(2, 121)    <= sub_wire6(121);
	sub_wire1(2, 122)    <= sub_wire6(122);
	sub_wire1(2, 123)    <= sub_wire6(123);
	sub_wire1(2, 124)    <= sub_wire6(124);
	sub_wire1(2, 125)    <= sub_wire6(125);
	sub_wire1(2, 126)    <= sub_wire6(126);
	sub_wire1(2, 127)    <= sub_wire6(127);
	sub_wire1(2, 128)    <= sub_wire6(128);
	sub_wire1(2, 129)    <= sub_wire6(129);
	sub_wire1(2, 130)    <= sub_wire6(130);
	sub_wire1(2, 131)    <= sub_wire6(131);
	sub_wire1(2, 132)    <= sub_wire6(132);
	sub_wire1(2, 133)    <= sub_wire6(133);
	sub_wire1(2, 134)    <= sub_wire6(134);
	sub_wire1(2, 135)    <= sub_wire6(135);
	sub_wire1(2, 136)    <= sub_wire6(136);
	sub_wire1(2, 137)    <= sub_wire6(137);
	sub_wire1(2, 138)    <= sub_wire6(138);
	sub_wire1(2, 139)    <= sub_wire6(139);
	sub_wire1(2, 140)    <= sub_wire6(140);
	sub_wire1(2, 141)    <= sub_wire6(141);
	sub_wire1(2, 142)    <= sub_wire6(142);
	sub_wire1(2, 143)    <= sub_wire6(143);
	sub_wire1(2, 144)    <= sub_wire6(144);
	sub_wire1(2, 145)    <= sub_wire6(145);
	sub_wire1(2, 146)    <= sub_wire6(146);
	sub_wire1(2, 147)    <= sub_wire6(147);
	sub_wire1(2, 148)    <= sub_wire6(148);
	sub_wire1(2, 149)    <= sub_wire6(149);
	sub_wire1(2, 150)    <= sub_wire6(150);
	sub_wire1(2, 151)    <= sub_wire6(151);
	sub_wire1(2, 152)    <= sub_wire6(152);
	sub_wire1(2, 153)    <= sub_wire6(153);
	sub_wire1(2, 154)    <= sub_wire6(154);
	sub_wire1(2, 155)    <= sub_wire6(155);
	sub_wire1(2, 156)    <= sub_wire6(156);
	sub_wire1(2, 157)    <= sub_wire6(157);
	sub_wire1(2, 158)    <= sub_wire6(158);
	sub_wire1(2, 159)    <= sub_wire6(159);
	sub_wire1(2, 160)    <= sub_wire6(160);
	sub_wire1(2, 161)    <= sub_wire6(161);
	sub_wire1(2, 162)    <= sub_wire6(162);
	sub_wire1(2, 163)    <= sub_wire6(163);
	sub_wire1(2, 164)    <= sub_wire6(164);
	sub_wire1(2, 165)    <= sub_wire6(165);
	sub_wire1(2, 166)    <= sub_wire6(166);
	sub_wire1(2, 167)    <= sub_wire6(167);
	sub_wire1(2, 168)    <= sub_wire6(168);
	sub_wire1(2, 169)    <= sub_wire6(169);
	sub_wire1(2, 170)    <= sub_wire6(170);
	sub_wire1(2, 171)    <= sub_wire6(171);
	sub_wire1(2, 172)    <= sub_wire6(172);
	sub_wire1(2, 173)    <= sub_wire6(173);
	sub_wire1(2, 174)    <= sub_wire6(174);
	sub_wire1(2, 175)    <= sub_wire6(175);
	sub_wire1(2, 176)    <= sub_wire6(176);
	sub_wire1(2, 177)    <= sub_wire6(177);
	sub_wire1(2, 178)    <= sub_wire6(178);
	sub_wire1(2, 179)    <= sub_wire6(179);
	sub_wire1(2, 180)    <= sub_wire6(180);
	sub_wire1(2, 181)    <= sub_wire6(181);
	sub_wire1(2, 182)    <= sub_wire6(182);
	sub_wire1(2, 183)    <= sub_wire6(183);
	sub_wire1(2, 184)    <= sub_wire6(184);
	sub_wire1(2, 185)    <= sub_wire6(185);
	sub_wire1(2, 186)    <= sub_wire6(186);
	sub_wire1(2, 187)    <= sub_wire6(187);
	sub_wire1(2, 188)    <= sub_wire6(188);
	sub_wire1(2, 189)    <= sub_wire6(189);
	sub_wire1(2, 190)    <= sub_wire6(190);
	sub_wire1(2, 191)    <= sub_wire6(191);
	sub_wire1(2, 192)    <= sub_wire6(192);
	sub_wire1(2, 193)    <= sub_wire6(193);
	sub_wire1(2, 194)    <= sub_wire6(194);
	sub_wire1(2, 195)    <= sub_wire6(195);
	sub_wire1(2, 196)    <= sub_wire6(196);
	sub_wire1(2, 197)    <= sub_wire6(197);
	sub_wire1(2, 198)    <= sub_wire6(198);
	sub_wire1(2, 199)    <= sub_wire6(199);
	sub_wire1(2, 200)    <= sub_wire6(200);
	sub_wire1(2, 201)    <= sub_wire6(201);
	sub_wire1(2, 202)    <= sub_wire6(202);
	sub_wire1(2, 203)    <= sub_wire6(203);
	sub_wire1(2, 204)    <= sub_wire6(204);
	sub_wire1(2, 205)    <= sub_wire6(205);
	sub_wire1(2, 206)    <= sub_wire6(206);
	sub_wire1(2, 207)    <= sub_wire6(207);
	sub_wire1(2, 208)    <= sub_wire6(208);
	sub_wire1(2, 209)    <= sub_wire6(209);
	sub_wire1(2, 210)    <= sub_wire6(210);
	sub_wire1(2, 211)    <= sub_wire6(211);
	sub_wire1(2, 212)    <= sub_wire6(212);
	sub_wire1(2, 213)    <= sub_wire6(213);
	sub_wire1(2, 214)    <= sub_wire6(214);
	sub_wire1(2, 215)    <= sub_wire6(215);
	sub_wire1(2, 216)    <= sub_wire6(216);
	sub_wire1(2, 217)    <= sub_wire6(217);
	sub_wire1(2, 218)    <= sub_wire6(218);
	sub_wire1(2, 219)    <= sub_wire6(219);
	sub_wire1(2, 220)    <= sub_wire6(220);
	sub_wire1(2, 221)    <= sub_wire6(221);
	sub_wire1(2, 222)    <= sub_wire6(222);
	sub_wire1(2, 223)    <= sub_wire6(223);
	sub_wire1(2, 224)    <= sub_wire6(224);
	sub_wire1(2, 225)    <= sub_wire6(225);
	sub_wire1(2, 226)    <= sub_wire6(226);
	sub_wire1(2, 227)    <= sub_wire6(227);
	sub_wire1(2, 228)    <= sub_wire6(228);
	sub_wire1(2, 229)    <= sub_wire6(229);
	sub_wire1(2, 230)    <= sub_wire6(230);
	sub_wire1(2, 231)    <= sub_wire6(231);
	sub_wire1(2, 232)    <= sub_wire6(232);
	sub_wire1(2, 233)    <= sub_wire6(233);
	sub_wire1(2, 234)    <= sub_wire6(234);
	sub_wire1(2, 235)    <= sub_wire6(235);
	sub_wire1(2, 236)    <= sub_wire6(236);
	sub_wire1(2, 237)    <= sub_wire6(237);
	sub_wire1(2, 238)    <= sub_wire6(238);
	sub_wire1(2, 239)    <= sub_wire6(239);
	sub_wire1(2, 240)    <= sub_wire6(240);
	sub_wire1(2, 241)    <= sub_wire6(241);
	sub_wire1(2, 242)    <= sub_wire6(242);
	sub_wire1(2, 243)    <= sub_wire6(243);
	sub_wire1(2, 244)    <= sub_wire6(244);
	sub_wire1(2, 245)    <= sub_wire6(245);
	sub_wire1(2, 246)    <= sub_wire6(246);
	sub_wire1(2, 247)    <= sub_wire6(247);
	sub_wire1(2, 248)    <= sub_wire6(248);
	sub_wire1(2, 249)    <= sub_wire6(249);
	sub_wire1(2, 250)    <= sub_wire6(250);
	sub_wire1(2, 251)    <= sub_wire6(251);
	sub_wire1(2, 252)    <= sub_wire6(252);
	sub_wire1(2, 253)    <= sub_wire6(253);
	sub_wire1(2, 254)    <= sub_wire6(254);
	sub_wire1(2, 255)    <= sub_wire6(255);
	sub_wire1(1, 0)    <= sub_wire7(0);
	sub_wire1(1, 1)    <= sub_wire7(1);
	sub_wire1(1, 2)    <= sub_wire7(2);
	sub_wire1(1, 3)    <= sub_wire7(3);
	sub_wire1(1, 4)    <= sub_wire7(4);
	sub_wire1(1, 5)    <= sub_wire7(5);
	sub_wire1(1, 6)    <= sub_wire7(6);
	sub_wire1(1, 7)    <= sub_wire7(7);
	sub_wire1(1, 8)    <= sub_wire7(8);
	sub_wire1(1, 9)    <= sub_wire7(9);
	sub_wire1(1, 10)    <= sub_wire7(10);
	sub_wire1(1, 11)    <= sub_wire7(11);
	sub_wire1(1, 12)    <= sub_wire7(12);
	sub_wire1(1, 13)    <= sub_wire7(13);
	sub_wire1(1, 14)    <= sub_wire7(14);
	sub_wire1(1, 15)    <= sub_wire7(15);
	sub_wire1(1, 16)    <= sub_wire7(16);
	sub_wire1(1, 17)    <= sub_wire7(17);
	sub_wire1(1, 18)    <= sub_wire7(18);
	sub_wire1(1, 19)    <= sub_wire7(19);
	sub_wire1(1, 20)    <= sub_wire7(20);
	sub_wire1(1, 21)    <= sub_wire7(21);
	sub_wire1(1, 22)    <= sub_wire7(22);
	sub_wire1(1, 23)    <= sub_wire7(23);
	sub_wire1(1, 24)    <= sub_wire7(24);
	sub_wire1(1, 25)    <= sub_wire7(25);
	sub_wire1(1, 26)    <= sub_wire7(26);
	sub_wire1(1, 27)    <= sub_wire7(27);
	sub_wire1(1, 28)    <= sub_wire7(28);
	sub_wire1(1, 29)    <= sub_wire7(29);
	sub_wire1(1, 30)    <= sub_wire7(30);
	sub_wire1(1, 31)    <= sub_wire7(31);
	sub_wire1(1, 32)    <= sub_wire7(32);
	sub_wire1(1, 33)    <= sub_wire7(33);
	sub_wire1(1, 34)    <= sub_wire7(34);
	sub_wire1(1, 35)    <= sub_wire7(35);
	sub_wire1(1, 36)    <= sub_wire7(36);
	sub_wire1(1, 37)    <= sub_wire7(37);
	sub_wire1(1, 38)    <= sub_wire7(38);
	sub_wire1(1, 39)    <= sub_wire7(39);
	sub_wire1(1, 40)    <= sub_wire7(40);
	sub_wire1(1, 41)    <= sub_wire7(41);
	sub_wire1(1, 42)    <= sub_wire7(42);
	sub_wire1(1, 43)    <= sub_wire7(43);
	sub_wire1(1, 44)    <= sub_wire7(44);
	sub_wire1(1, 45)    <= sub_wire7(45);
	sub_wire1(1, 46)    <= sub_wire7(46);
	sub_wire1(1, 47)    <= sub_wire7(47);
	sub_wire1(1, 48)    <= sub_wire7(48);
	sub_wire1(1, 49)    <= sub_wire7(49);
	sub_wire1(1, 50)    <= sub_wire7(50);
	sub_wire1(1, 51)    <= sub_wire7(51);
	sub_wire1(1, 52)    <= sub_wire7(52);
	sub_wire1(1, 53)    <= sub_wire7(53);
	sub_wire1(1, 54)    <= sub_wire7(54);
	sub_wire1(1, 55)    <= sub_wire7(55);
	sub_wire1(1, 56)    <= sub_wire7(56);
	sub_wire1(1, 57)    <= sub_wire7(57);
	sub_wire1(1, 58)    <= sub_wire7(58);
	sub_wire1(1, 59)    <= sub_wire7(59);
	sub_wire1(1, 60)    <= sub_wire7(60);
	sub_wire1(1, 61)    <= sub_wire7(61);
	sub_wire1(1, 62)    <= sub_wire7(62);
	sub_wire1(1, 63)    <= sub_wire7(63);
	sub_wire1(1, 64)    <= sub_wire7(64);
	sub_wire1(1, 65)    <= sub_wire7(65);
	sub_wire1(1, 66)    <= sub_wire7(66);
	sub_wire1(1, 67)    <= sub_wire7(67);
	sub_wire1(1, 68)    <= sub_wire7(68);
	sub_wire1(1, 69)    <= sub_wire7(69);
	sub_wire1(1, 70)    <= sub_wire7(70);
	sub_wire1(1, 71)    <= sub_wire7(71);
	sub_wire1(1, 72)    <= sub_wire7(72);
	sub_wire1(1, 73)    <= sub_wire7(73);
	sub_wire1(1, 74)    <= sub_wire7(74);
	sub_wire1(1, 75)    <= sub_wire7(75);
	sub_wire1(1, 76)    <= sub_wire7(76);
	sub_wire1(1, 77)    <= sub_wire7(77);
	sub_wire1(1, 78)    <= sub_wire7(78);
	sub_wire1(1, 79)    <= sub_wire7(79);
	sub_wire1(1, 80)    <= sub_wire7(80);
	sub_wire1(1, 81)    <= sub_wire7(81);
	sub_wire1(1, 82)    <= sub_wire7(82);
	sub_wire1(1, 83)    <= sub_wire7(83);
	sub_wire1(1, 84)    <= sub_wire7(84);
	sub_wire1(1, 85)    <= sub_wire7(85);
	sub_wire1(1, 86)    <= sub_wire7(86);
	sub_wire1(1, 87)    <= sub_wire7(87);
	sub_wire1(1, 88)    <= sub_wire7(88);
	sub_wire1(1, 89)    <= sub_wire7(89);
	sub_wire1(1, 90)    <= sub_wire7(90);
	sub_wire1(1, 91)    <= sub_wire7(91);
	sub_wire1(1, 92)    <= sub_wire7(92);
	sub_wire1(1, 93)    <= sub_wire7(93);
	sub_wire1(1, 94)    <= sub_wire7(94);
	sub_wire1(1, 95)    <= sub_wire7(95);
	sub_wire1(1, 96)    <= sub_wire7(96);
	sub_wire1(1, 97)    <= sub_wire7(97);
	sub_wire1(1, 98)    <= sub_wire7(98);
	sub_wire1(1, 99)    <= sub_wire7(99);
	sub_wire1(1, 100)    <= sub_wire7(100);
	sub_wire1(1, 101)    <= sub_wire7(101);
	sub_wire1(1, 102)    <= sub_wire7(102);
	sub_wire1(1, 103)    <= sub_wire7(103);
	sub_wire1(1, 104)    <= sub_wire7(104);
	sub_wire1(1, 105)    <= sub_wire7(105);
	sub_wire1(1, 106)    <= sub_wire7(106);
	sub_wire1(1, 107)    <= sub_wire7(107);
	sub_wire1(1, 108)    <= sub_wire7(108);
	sub_wire1(1, 109)    <= sub_wire7(109);
	sub_wire1(1, 110)    <= sub_wire7(110);
	sub_wire1(1, 111)    <= sub_wire7(111);
	sub_wire1(1, 112)    <= sub_wire7(112);
	sub_wire1(1, 113)    <= sub_wire7(113);
	sub_wire1(1, 114)    <= sub_wire7(114);
	sub_wire1(1, 115)    <= sub_wire7(115);
	sub_wire1(1, 116)    <= sub_wire7(116);
	sub_wire1(1, 117)    <= sub_wire7(117);
	sub_wire1(1, 118)    <= sub_wire7(118);
	sub_wire1(1, 119)    <= sub_wire7(119);
	sub_wire1(1, 120)    <= sub_wire7(120);
	sub_wire1(1, 121)    <= sub_wire7(121);
	sub_wire1(1, 122)    <= sub_wire7(122);
	sub_wire1(1, 123)    <= sub_wire7(123);
	sub_wire1(1, 124)    <= sub_wire7(124);
	sub_wire1(1, 125)    <= sub_wire7(125);
	sub_wire1(1, 126)    <= sub_wire7(126);
	sub_wire1(1, 127)    <= sub_wire7(127);
	sub_wire1(1, 128)    <= sub_wire7(128);
	sub_wire1(1, 129)    <= sub_wire7(129);
	sub_wire1(1, 130)    <= sub_wire7(130);
	sub_wire1(1, 131)    <= sub_wire7(131);
	sub_wire1(1, 132)    <= sub_wire7(132);
	sub_wire1(1, 133)    <= sub_wire7(133);
	sub_wire1(1, 134)    <= sub_wire7(134);
	sub_wire1(1, 135)    <= sub_wire7(135);
	sub_wire1(1, 136)    <= sub_wire7(136);
	sub_wire1(1, 137)    <= sub_wire7(137);
	sub_wire1(1, 138)    <= sub_wire7(138);
	sub_wire1(1, 139)    <= sub_wire7(139);
	sub_wire1(1, 140)    <= sub_wire7(140);
	sub_wire1(1, 141)    <= sub_wire7(141);
	sub_wire1(1, 142)    <= sub_wire7(142);
	sub_wire1(1, 143)    <= sub_wire7(143);
	sub_wire1(1, 144)    <= sub_wire7(144);
	sub_wire1(1, 145)    <= sub_wire7(145);
	sub_wire1(1, 146)    <= sub_wire7(146);
	sub_wire1(1, 147)    <= sub_wire7(147);
	sub_wire1(1, 148)    <= sub_wire7(148);
	sub_wire1(1, 149)    <= sub_wire7(149);
	sub_wire1(1, 150)    <= sub_wire7(150);
	sub_wire1(1, 151)    <= sub_wire7(151);
	sub_wire1(1, 152)    <= sub_wire7(152);
	sub_wire1(1, 153)    <= sub_wire7(153);
	sub_wire1(1, 154)    <= sub_wire7(154);
	sub_wire1(1, 155)    <= sub_wire7(155);
	sub_wire1(1, 156)    <= sub_wire7(156);
	sub_wire1(1, 157)    <= sub_wire7(157);
	sub_wire1(1, 158)    <= sub_wire7(158);
	sub_wire1(1, 159)    <= sub_wire7(159);
	sub_wire1(1, 160)    <= sub_wire7(160);
	sub_wire1(1, 161)    <= sub_wire7(161);
	sub_wire1(1, 162)    <= sub_wire7(162);
	sub_wire1(1, 163)    <= sub_wire7(163);
	sub_wire1(1, 164)    <= sub_wire7(164);
	sub_wire1(1, 165)    <= sub_wire7(165);
	sub_wire1(1, 166)    <= sub_wire7(166);
	sub_wire1(1, 167)    <= sub_wire7(167);
	sub_wire1(1, 168)    <= sub_wire7(168);
	sub_wire1(1, 169)    <= sub_wire7(169);
	sub_wire1(1, 170)    <= sub_wire7(170);
	sub_wire1(1, 171)    <= sub_wire7(171);
	sub_wire1(1, 172)    <= sub_wire7(172);
	sub_wire1(1, 173)    <= sub_wire7(173);
	sub_wire1(1, 174)    <= sub_wire7(174);
	sub_wire1(1, 175)    <= sub_wire7(175);
	sub_wire1(1, 176)    <= sub_wire7(176);
	sub_wire1(1, 177)    <= sub_wire7(177);
	sub_wire1(1, 178)    <= sub_wire7(178);
	sub_wire1(1, 179)    <= sub_wire7(179);
	sub_wire1(1, 180)    <= sub_wire7(180);
	sub_wire1(1, 181)    <= sub_wire7(181);
	sub_wire1(1, 182)    <= sub_wire7(182);
	sub_wire1(1, 183)    <= sub_wire7(183);
	sub_wire1(1, 184)    <= sub_wire7(184);
	sub_wire1(1, 185)    <= sub_wire7(185);
	sub_wire1(1, 186)    <= sub_wire7(186);
	sub_wire1(1, 187)    <= sub_wire7(187);
	sub_wire1(1, 188)    <= sub_wire7(188);
	sub_wire1(1, 189)    <= sub_wire7(189);
	sub_wire1(1, 190)    <= sub_wire7(190);
	sub_wire1(1, 191)    <= sub_wire7(191);
	sub_wire1(1, 192)    <= sub_wire7(192);
	sub_wire1(1, 193)    <= sub_wire7(193);
	sub_wire1(1, 194)    <= sub_wire7(194);
	sub_wire1(1, 195)    <= sub_wire7(195);
	sub_wire1(1, 196)    <= sub_wire7(196);
	sub_wire1(1, 197)    <= sub_wire7(197);
	sub_wire1(1, 198)    <= sub_wire7(198);
	sub_wire1(1, 199)    <= sub_wire7(199);
	sub_wire1(1, 200)    <= sub_wire7(200);
	sub_wire1(1, 201)    <= sub_wire7(201);
	sub_wire1(1, 202)    <= sub_wire7(202);
	sub_wire1(1, 203)    <= sub_wire7(203);
	sub_wire1(1, 204)    <= sub_wire7(204);
	sub_wire1(1, 205)    <= sub_wire7(205);
	sub_wire1(1, 206)    <= sub_wire7(206);
	sub_wire1(1, 207)    <= sub_wire7(207);
	sub_wire1(1, 208)    <= sub_wire7(208);
	sub_wire1(1, 209)    <= sub_wire7(209);
	sub_wire1(1, 210)    <= sub_wire7(210);
	sub_wire1(1, 211)    <= sub_wire7(211);
	sub_wire1(1, 212)    <= sub_wire7(212);
	sub_wire1(1, 213)    <= sub_wire7(213);
	sub_wire1(1, 214)    <= sub_wire7(214);
	sub_wire1(1, 215)    <= sub_wire7(215);
	sub_wire1(1, 216)    <= sub_wire7(216);
	sub_wire1(1, 217)    <= sub_wire7(217);
	sub_wire1(1, 218)    <= sub_wire7(218);
	sub_wire1(1, 219)    <= sub_wire7(219);
	sub_wire1(1, 220)    <= sub_wire7(220);
	sub_wire1(1, 221)    <= sub_wire7(221);
	sub_wire1(1, 222)    <= sub_wire7(222);
	sub_wire1(1, 223)    <= sub_wire7(223);
	sub_wire1(1, 224)    <= sub_wire7(224);
	sub_wire1(1, 225)    <= sub_wire7(225);
	sub_wire1(1, 226)    <= sub_wire7(226);
	sub_wire1(1, 227)    <= sub_wire7(227);
	sub_wire1(1, 228)    <= sub_wire7(228);
	sub_wire1(1, 229)    <= sub_wire7(229);
	sub_wire1(1, 230)    <= sub_wire7(230);
	sub_wire1(1, 231)    <= sub_wire7(231);
	sub_wire1(1, 232)    <= sub_wire7(232);
	sub_wire1(1, 233)    <= sub_wire7(233);
	sub_wire1(1, 234)    <= sub_wire7(234);
	sub_wire1(1, 235)    <= sub_wire7(235);
	sub_wire1(1, 236)    <= sub_wire7(236);
	sub_wire1(1, 237)    <= sub_wire7(237);
	sub_wire1(1, 238)    <= sub_wire7(238);
	sub_wire1(1, 239)    <= sub_wire7(239);
	sub_wire1(1, 240)    <= sub_wire7(240);
	sub_wire1(1, 241)    <= sub_wire7(241);
	sub_wire1(1, 242)    <= sub_wire7(242);
	sub_wire1(1, 243)    <= sub_wire7(243);
	sub_wire1(1, 244)    <= sub_wire7(244);
	sub_wire1(1, 245)    <= sub_wire7(245);
	sub_wire1(1, 246)    <= sub_wire7(246);
	sub_wire1(1, 247)    <= sub_wire7(247);
	sub_wire1(1, 248)    <= sub_wire7(248);
	sub_wire1(1, 249)    <= sub_wire7(249);
	sub_wire1(1, 250)    <= sub_wire7(250);
	sub_wire1(1, 251)    <= sub_wire7(251);
	sub_wire1(1, 252)    <= sub_wire7(252);
	sub_wire1(1, 253)    <= sub_wire7(253);
	sub_wire1(1, 254)    <= sub_wire7(254);
	sub_wire1(1, 255)    <= sub_wire7(255);
	sub_wire1(0, 0)    <= sub_wire8(0);
	sub_wire1(0, 1)    <= sub_wire8(1);
	sub_wire1(0, 2)    <= sub_wire8(2);
	sub_wire1(0, 3)    <= sub_wire8(3);
	sub_wire1(0, 4)    <= sub_wire8(4);
	sub_wire1(0, 5)    <= sub_wire8(5);
	sub_wire1(0, 6)    <= sub_wire8(6);
	sub_wire1(0, 7)    <= sub_wire8(7);
	sub_wire1(0, 8)    <= sub_wire8(8);
	sub_wire1(0, 9)    <= sub_wire8(9);
	sub_wire1(0, 10)    <= sub_wire8(10);
	sub_wire1(0, 11)    <= sub_wire8(11);
	sub_wire1(0, 12)    <= sub_wire8(12);
	sub_wire1(0, 13)    <= sub_wire8(13);
	sub_wire1(0, 14)    <= sub_wire8(14);
	sub_wire1(0, 15)    <= sub_wire8(15);
	sub_wire1(0, 16)    <= sub_wire8(16);
	sub_wire1(0, 17)    <= sub_wire8(17);
	sub_wire1(0, 18)    <= sub_wire8(18);
	sub_wire1(0, 19)    <= sub_wire8(19);
	sub_wire1(0, 20)    <= sub_wire8(20);
	sub_wire1(0, 21)    <= sub_wire8(21);
	sub_wire1(0, 22)    <= sub_wire8(22);
	sub_wire1(0, 23)    <= sub_wire8(23);
	sub_wire1(0, 24)    <= sub_wire8(24);
	sub_wire1(0, 25)    <= sub_wire8(25);
	sub_wire1(0, 26)    <= sub_wire8(26);
	sub_wire1(0, 27)    <= sub_wire8(27);
	sub_wire1(0, 28)    <= sub_wire8(28);
	sub_wire1(0, 29)    <= sub_wire8(29);
	sub_wire1(0, 30)    <= sub_wire8(30);
	sub_wire1(0, 31)    <= sub_wire8(31);
	sub_wire1(0, 32)    <= sub_wire8(32);
	sub_wire1(0, 33)    <= sub_wire8(33);
	sub_wire1(0, 34)    <= sub_wire8(34);
	sub_wire1(0, 35)    <= sub_wire8(35);
	sub_wire1(0, 36)    <= sub_wire8(36);
	sub_wire1(0, 37)    <= sub_wire8(37);
	sub_wire1(0, 38)    <= sub_wire8(38);
	sub_wire1(0, 39)    <= sub_wire8(39);
	sub_wire1(0, 40)    <= sub_wire8(40);
	sub_wire1(0, 41)    <= sub_wire8(41);
	sub_wire1(0, 42)    <= sub_wire8(42);
	sub_wire1(0, 43)    <= sub_wire8(43);
	sub_wire1(0, 44)    <= sub_wire8(44);
	sub_wire1(0, 45)    <= sub_wire8(45);
	sub_wire1(0, 46)    <= sub_wire8(46);
	sub_wire1(0, 47)    <= sub_wire8(47);
	sub_wire1(0, 48)    <= sub_wire8(48);
	sub_wire1(0, 49)    <= sub_wire8(49);
	sub_wire1(0, 50)    <= sub_wire8(50);
	sub_wire1(0, 51)    <= sub_wire8(51);
	sub_wire1(0, 52)    <= sub_wire8(52);
	sub_wire1(0, 53)    <= sub_wire8(53);
	sub_wire1(0, 54)    <= sub_wire8(54);
	sub_wire1(0, 55)    <= sub_wire8(55);
	sub_wire1(0, 56)    <= sub_wire8(56);
	sub_wire1(0, 57)    <= sub_wire8(57);
	sub_wire1(0, 58)    <= sub_wire8(58);
	sub_wire1(0, 59)    <= sub_wire8(59);
	sub_wire1(0, 60)    <= sub_wire8(60);
	sub_wire1(0, 61)    <= sub_wire8(61);
	sub_wire1(0, 62)    <= sub_wire8(62);
	sub_wire1(0, 63)    <= sub_wire8(63);
	sub_wire1(0, 64)    <= sub_wire8(64);
	sub_wire1(0, 65)    <= sub_wire8(65);
	sub_wire1(0, 66)    <= sub_wire8(66);
	sub_wire1(0, 67)    <= sub_wire8(67);
	sub_wire1(0, 68)    <= sub_wire8(68);
	sub_wire1(0, 69)    <= sub_wire8(69);
	sub_wire1(0, 70)    <= sub_wire8(70);
	sub_wire1(0, 71)    <= sub_wire8(71);
	sub_wire1(0, 72)    <= sub_wire8(72);
	sub_wire1(0, 73)    <= sub_wire8(73);
	sub_wire1(0, 74)    <= sub_wire8(74);
	sub_wire1(0, 75)    <= sub_wire8(75);
	sub_wire1(0, 76)    <= sub_wire8(76);
	sub_wire1(0, 77)    <= sub_wire8(77);
	sub_wire1(0, 78)    <= sub_wire8(78);
	sub_wire1(0, 79)    <= sub_wire8(79);
	sub_wire1(0, 80)    <= sub_wire8(80);
	sub_wire1(0, 81)    <= sub_wire8(81);
	sub_wire1(0, 82)    <= sub_wire8(82);
	sub_wire1(0, 83)    <= sub_wire8(83);
	sub_wire1(0, 84)    <= sub_wire8(84);
	sub_wire1(0, 85)    <= sub_wire8(85);
	sub_wire1(0, 86)    <= sub_wire8(86);
	sub_wire1(0, 87)    <= sub_wire8(87);
	sub_wire1(0, 88)    <= sub_wire8(88);
	sub_wire1(0, 89)    <= sub_wire8(89);
	sub_wire1(0, 90)    <= sub_wire8(90);
	sub_wire1(0, 91)    <= sub_wire8(91);
	sub_wire1(0, 92)    <= sub_wire8(92);
	sub_wire1(0, 93)    <= sub_wire8(93);
	sub_wire1(0, 94)    <= sub_wire8(94);
	sub_wire1(0, 95)    <= sub_wire8(95);
	sub_wire1(0, 96)    <= sub_wire8(96);
	sub_wire1(0, 97)    <= sub_wire8(97);
	sub_wire1(0, 98)    <= sub_wire8(98);
	sub_wire1(0, 99)    <= sub_wire8(99);
	sub_wire1(0, 100)    <= sub_wire8(100);
	sub_wire1(0, 101)    <= sub_wire8(101);
	sub_wire1(0, 102)    <= sub_wire8(102);
	sub_wire1(0, 103)    <= sub_wire8(103);
	sub_wire1(0, 104)    <= sub_wire8(104);
	sub_wire1(0, 105)    <= sub_wire8(105);
	sub_wire1(0, 106)    <= sub_wire8(106);
	sub_wire1(0, 107)    <= sub_wire8(107);
	sub_wire1(0, 108)    <= sub_wire8(108);
	sub_wire1(0, 109)    <= sub_wire8(109);
	sub_wire1(0, 110)    <= sub_wire8(110);
	sub_wire1(0, 111)    <= sub_wire8(111);
	sub_wire1(0, 112)    <= sub_wire8(112);
	sub_wire1(0, 113)    <= sub_wire8(113);
	sub_wire1(0, 114)    <= sub_wire8(114);
	sub_wire1(0, 115)    <= sub_wire8(115);
	sub_wire1(0, 116)    <= sub_wire8(116);
	sub_wire1(0, 117)    <= sub_wire8(117);
	sub_wire1(0, 118)    <= sub_wire8(118);
	sub_wire1(0, 119)    <= sub_wire8(119);
	sub_wire1(0, 120)    <= sub_wire8(120);
	sub_wire1(0, 121)    <= sub_wire8(121);
	sub_wire1(0, 122)    <= sub_wire8(122);
	sub_wire1(0, 123)    <= sub_wire8(123);
	sub_wire1(0, 124)    <= sub_wire8(124);
	sub_wire1(0, 125)    <= sub_wire8(125);
	sub_wire1(0, 126)    <= sub_wire8(126);
	sub_wire1(0, 127)    <= sub_wire8(127);
	sub_wire1(0, 128)    <= sub_wire8(128);
	sub_wire1(0, 129)    <= sub_wire8(129);
	sub_wire1(0, 130)    <= sub_wire8(130);
	sub_wire1(0, 131)    <= sub_wire8(131);
	sub_wire1(0, 132)    <= sub_wire8(132);
	sub_wire1(0, 133)    <= sub_wire8(133);
	sub_wire1(0, 134)    <= sub_wire8(134);
	sub_wire1(0, 135)    <= sub_wire8(135);
	sub_wire1(0, 136)    <= sub_wire8(136);
	sub_wire1(0, 137)    <= sub_wire8(137);
	sub_wire1(0, 138)    <= sub_wire8(138);
	sub_wire1(0, 139)    <= sub_wire8(139);
	sub_wire1(0, 140)    <= sub_wire8(140);
	sub_wire1(0, 141)    <= sub_wire8(141);
	sub_wire1(0, 142)    <= sub_wire8(142);
	sub_wire1(0, 143)    <= sub_wire8(143);
	sub_wire1(0, 144)    <= sub_wire8(144);
	sub_wire1(0, 145)    <= sub_wire8(145);
	sub_wire1(0, 146)    <= sub_wire8(146);
	sub_wire1(0, 147)    <= sub_wire8(147);
	sub_wire1(0, 148)    <= sub_wire8(148);
	sub_wire1(0, 149)    <= sub_wire8(149);
	sub_wire1(0, 150)    <= sub_wire8(150);
	sub_wire1(0, 151)    <= sub_wire8(151);
	sub_wire1(0, 152)    <= sub_wire8(152);
	sub_wire1(0, 153)    <= sub_wire8(153);
	sub_wire1(0, 154)    <= sub_wire8(154);
	sub_wire1(0, 155)    <= sub_wire8(155);
	sub_wire1(0, 156)    <= sub_wire8(156);
	sub_wire1(0, 157)    <= sub_wire8(157);
	sub_wire1(0, 158)    <= sub_wire8(158);
	sub_wire1(0, 159)    <= sub_wire8(159);
	sub_wire1(0, 160)    <= sub_wire8(160);
	sub_wire1(0, 161)    <= sub_wire8(161);
	sub_wire1(0, 162)    <= sub_wire8(162);
	sub_wire1(0, 163)    <= sub_wire8(163);
	sub_wire1(0, 164)    <= sub_wire8(164);
	sub_wire1(0, 165)    <= sub_wire8(165);
	sub_wire1(0, 166)    <= sub_wire8(166);
	sub_wire1(0, 167)    <= sub_wire8(167);
	sub_wire1(0, 168)    <= sub_wire8(168);
	sub_wire1(0, 169)    <= sub_wire8(169);
	sub_wire1(0, 170)    <= sub_wire8(170);
	sub_wire1(0, 171)    <= sub_wire8(171);
	sub_wire1(0, 172)    <= sub_wire8(172);
	sub_wire1(0, 173)    <= sub_wire8(173);
	sub_wire1(0, 174)    <= sub_wire8(174);
	sub_wire1(0, 175)    <= sub_wire8(175);
	sub_wire1(0, 176)    <= sub_wire8(176);
	sub_wire1(0, 177)    <= sub_wire8(177);
	sub_wire1(0, 178)    <= sub_wire8(178);
	sub_wire1(0, 179)    <= sub_wire8(179);
	sub_wire1(0, 180)    <= sub_wire8(180);
	sub_wire1(0, 181)    <= sub_wire8(181);
	sub_wire1(0, 182)    <= sub_wire8(182);
	sub_wire1(0, 183)    <= sub_wire8(183);
	sub_wire1(0, 184)    <= sub_wire8(184);
	sub_wire1(0, 185)    <= sub_wire8(185);
	sub_wire1(0, 186)    <= sub_wire8(186);
	sub_wire1(0, 187)    <= sub_wire8(187);
	sub_wire1(0, 188)    <= sub_wire8(188);
	sub_wire1(0, 189)    <= sub_wire8(189);
	sub_wire1(0, 190)    <= sub_wire8(190);
	sub_wire1(0, 191)    <= sub_wire8(191);
	sub_wire1(0, 192)    <= sub_wire8(192);
	sub_wire1(0, 193)    <= sub_wire8(193);
	sub_wire1(0, 194)    <= sub_wire8(194);
	sub_wire1(0, 195)    <= sub_wire8(195);
	sub_wire1(0, 196)    <= sub_wire8(196);
	sub_wire1(0, 197)    <= sub_wire8(197);
	sub_wire1(0, 198)    <= sub_wire8(198);
	sub_wire1(0, 199)    <= sub_wire8(199);
	sub_wire1(0, 200)    <= sub_wire8(200);
	sub_wire1(0, 201)    <= sub_wire8(201);
	sub_wire1(0, 202)    <= sub_wire8(202);
	sub_wire1(0, 203)    <= sub_wire8(203);
	sub_wire1(0, 204)    <= sub_wire8(204);
	sub_wire1(0, 205)    <= sub_wire8(205);
	sub_wire1(0, 206)    <= sub_wire8(206);
	sub_wire1(0, 207)    <= sub_wire8(207);
	sub_wire1(0, 208)    <= sub_wire8(208);
	sub_wire1(0, 209)    <= sub_wire8(209);
	sub_wire1(0, 210)    <= sub_wire8(210);
	sub_wire1(0, 211)    <= sub_wire8(211);
	sub_wire1(0, 212)    <= sub_wire8(212);
	sub_wire1(0, 213)    <= sub_wire8(213);
	sub_wire1(0, 214)    <= sub_wire8(214);
	sub_wire1(0, 215)    <= sub_wire8(215);
	sub_wire1(0, 216)    <= sub_wire8(216);
	sub_wire1(0, 217)    <= sub_wire8(217);
	sub_wire1(0, 218)    <= sub_wire8(218);
	sub_wire1(0, 219)    <= sub_wire8(219);
	sub_wire1(0, 220)    <= sub_wire8(220);
	sub_wire1(0, 221)    <= sub_wire8(221);
	sub_wire1(0, 222)    <= sub_wire8(222);
	sub_wire1(0, 223)    <= sub_wire8(223);
	sub_wire1(0, 224)    <= sub_wire8(224);
	sub_wire1(0, 225)    <= sub_wire8(225);
	sub_wire1(0, 226)    <= sub_wire8(226);
	sub_wire1(0, 227)    <= sub_wire8(227);
	sub_wire1(0, 228)    <= sub_wire8(228);
	sub_wire1(0, 229)    <= sub_wire8(229);
	sub_wire1(0, 230)    <= sub_wire8(230);
	sub_wire1(0, 231)    <= sub_wire8(231);
	sub_wire1(0, 232)    <= sub_wire8(232);
	sub_wire1(0, 233)    <= sub_wire8(233);
	sub_wire1(0, 234)    <= sub_wire8(234);
	sub_wire1(0, 235)    <= sub_wire8(235);
	sub_wire1(0, 236)    <= sub_wire8(236);
	sub_wire1(0, 237)    <= sub_wire8(237);
	sub_wire1(0, 238)    <= sub_wire8(238);
	sub_wire1(0, 239)    <= sub_wire8(239);
	sub_wire1(0, 240)    <= sub_wire8(240);
	sub_wire1(0, 241)    <= sub_wire8(241);
	sub_wire1(0, 242)    <= sub_wire8(242);
	sub_wire1(0, 243)    <= sub_wire8(243);
	sub_wire1(0, 244)    <= sub_wire8(244);
	sub_wire1(0, 245)    <= sub_wire8(245);
	sub_wire1(0, 246)    <= sub_wire8(246);
	sub_wire1(0, 247)    <= sub_wire8(247);
	sub_wire1(0, 248)    <= sub_wire8(248);
	sub_wire1(0, 249)    <= sub_wire8(249);
	sub_wire1(0, 250)    <= sub_wire8(250);
	sub_wire1(0, 251)    <= sub_wire8(251);
	sub_wire1(0, 252)    <= sub_wire8(252);
	sub_wire1(0, 253)    <= sub_wire8(253);
	sub_wire1(0, 254)    <= sub_wire8(254);
	sub_wire1(0, 255)    <= sub_wire8(255);
	result    <= sub_wire9(255 DOWNTO 0);

	LPM_MUX_component : LPM_MUX
	GENERIC MAP (
		lpm_pipeline => 1,
		lpm_size => 8,
		lpm_type => "LPM_MUX",
		lpm_width => 256,
		lpm_widths => 3
	)
	PORT MAP (
		clock => clock,
		data => sub_wire1,
		sel => sel,
		result => sub_wire9
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "1"
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "8"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "256"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "3"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data0x 0 0 256 0 INPUT NODEFVAL "data0x[255..0]"
-- Retrieval info: USED_PORT: data1x 0 0 256 0 INPUT NODEFVAL "data1x[255..0]"
-- Retrieval info: USED_PORT: data2x 0 0 256 0 INPUT NODEFVAL "data2x[255..0]"
-- Retrieval info: USED_PORT: data3x 0 0 256 0 INPUT NODEFVAL "data3x[255..0]"
-- Retrieval info: USED_PORT: data4x 0 0 256 0 INPUT NODEFVAL "data4x[255..0]"
-- Retrieval info: USED_PORT: data5x 0 0 256 0 INPUT NODEFVAL "data5x[255..0]"
-- Retrieval info: USED_PORT: data6x 0 0 256 0 INPUT NODEFVAL "data6x[255..0]"
-- Retrieval info: USED_PORT: data7x 0 0 256 0 INPUT NODEFVAL "data7x[255..0]"
-- Retrieval info: USED_PORT: result 0 0 256 0 OUTPUT NODEFVAL "result[255..0]"
-- Retrieval info: USED_PORT: sel 0 0 3 0 INPUT NODEFVAL "sel[2..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data 1 0 256 0 data0x 0 0 256 0
-- Retrieval info: CONNECT: @data 1 1 256 0 data1x 0 0 256 0
-- Retrieval info: CONNECT: @data 1 2 256 0 data2x 0 0 256 0
-- Retrieval info: CONNECT: @data 1 3 256 0 data3x 0 0 256 0
-- Retrieval info: CONNECT: @data 1 4 256 0 data4x 0 0 256 0
-- Retrieval info: CONNECT: @data 1 5 256 0 data5x 0 0 256 0
-- Retrieval info: CONNECT: @data 1 6 256 0 data6x 0 0 256 0
-- Retrieval info: CONNECT: @data 1 7 256 0 data7x 0 0 256 0
-- Retrieval info: CONNECT: @sel 0 0 3 0 sel 0 0 3 0
-- Retrieval info: CONNECT: result 0 0 256 0 @result 0 0 256 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX8_256b.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX8_256b.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX8_256b.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX8_256b.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX8_256b_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
