-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_MUX 

-- ============================================================
-- File Name: mux256.vhd
-- Megafunction Name(s):
-- 			LPM_MUX
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.0 Build 156 04/24/2013 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY mux256 IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		sel		: IN STD_LOGIC ;
		result		: OUT STD_LOGIC_VECTOR (255 DOWNTO 0)
	);
END mux256;


ARCHITECTURE SYN OF mux256 IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_2D (1 DOWNTO 0, 255 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (255 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC ;
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (0 DOWNTO 0);

BEGIN
	sub_wire3    <= data0x(255 DOWNTO 0);
	result    <= sub_wire0(255 DOWNTO 0);
	sub_wire1    <= data1x(255 DOWNTO 0);
	sub_wire2(1, 0)    <= sub_wire1(0);
	sub_wire2(1, 1)    <= sub_wire1(1);
	sub_wire2(1, 2)    <= sub_wire1(2);
	sub_wire2(1, 3)    <= sub_wire1(3);
	sub_wire2(1, 4)    <= sub_wire1(4);
	sub_wire2(1, 5)    <= sub_wire1(5);
	sub_wire2(1, 6)    <= sub_wire1(6);
	sub_wire2(1, 7)    <= sub_wire1(7);
	sub_wire2(1, 8)    <= sub_wire1(8);
	sub_wire2(1, 9)    <= sub_wire1(9);
	sub_wire2(1, 10)    <= sub_wire1(10);
	sub_wire2(1, 11)    <= sub_wire1(11);
	sub_wire2(1, 12)    <= sub_wire1(12);
	sub_wire2(1, 13)    <= sub_wire1(13);
	sub_wire2(1, 14)    <= sub_wire1(14);
	sub_wire2(1, 15)    <= sub_wire1(15);
	sub_wire2(1, 16)    <= sub_wire1(16);
	sub_wire2(1, 17)    <= sub_wire1(17);
	sub_wire2(1, 18)    <= sub_wire1(18);
	sub_wire2(1, 19)    <= sub_wire1(19);
	sub_wire2(1, 20)    <= sub_wire1(20);
	sub_wire2(1, 21)    <= sub_wire1(21);
	sub_wire2(1, 22)    <= sub_wire1(22);
	sub_wire2(1, 23)    <= sub_wire1(23);
	sub_wire2(1, 24)    <= sub_wire1(24);
	sub_wire2(1, 25)    <= sub_wire1(25);
	sub_wire2(1, 26)    <= sub_wire1(26);
	sub_wire2(1, 27)    <= sub_wire1(27);
	sub_wire2(1, 28)    <= sub_wire1(28);
	sub_wire2(1, 29)    <= sub_wire1(29);
	sub_wire2(1, 30)    <= sub_wire1(30);
	sub_wire2(1, 31)    <= sub_wire1(31);
	sub_wire2(1, 32)    <= sub_wire1(32);
	sub_wire2(1, 33)    <= sub_wire1(33);
	sub_wire2(1, 34)    <= sub_wire1(34);
	sub_wire2(1, 35)    <= sub_wire1(35);
	sub_wire2(1, 36)    <= sub_wire1(36);
	sub_wire2(1, 37)    <= sub_wire1(37);
	sub_wire2(1, 38)    <= sub_wire1(38);
	sub_wire2(1, 39)    <= sub_wire1(39);
	sub_wire2(1, 40)    <= sub_wire1(40);
	sub_wire2(1, 41)    <= sub_wire1(41);
	sub_wire2(1, 42)    <= sub_wire1(42);
	sub_wire2(1, 43)    <= sub_wire1(43);
	sub_wire2(1, 44)    <= sub_wire1(44);
	sub_wire2(1, 45)    <= sub_wire1(45);
	sub_wire2(1, 46)    <= sub_wire1(46);
	sub_wire2(1, 47)    <= sub_wire1(47);
	sub_wire2(1, 48)    <= sub_wire1(48);
	sub_wire2(1, 49)    <= sub_wire1(49);
	sub_wire2(1, 50)    <= sub_wire1(50);
	sub_wire2(1, 51)    <= sub_wire1(51);
	sub_wire2(1, 52)    <= sub_wire1(52);
	sub_wire2(1, 53)    <= sub_wire1(53);
	sub_wire2(1, 54)    <= sub_wire1(54);
	sub_wire2(1, 55)    <= sub_wire1(55);
	sub_wire2(1, 56)    <= sub_wire1(56);
	sub_wire2(1, 57)    <= sub_wire1(57);
	sub_wire2(1, 58)    <= sub_wire1(58);
	sub_wire2(1, 59)    <= sub_wire1(59);
	sub_wire2(1, 60)    <= sub_wire1(60);
	sub_wire2(1, 61)    <= sub_wire1(61);
	sub_wire2(1, 62)    <= sub_wire1(62);
	sub_wire2(1, 63)    <= sub_wire1(63);
	sub_wire2(1, 64)    <= sub_wire1(64);
	sub_wire2(1, 65)    <= sub_wire1(65);
	sub_wire2(1, 66)    <= sub_wire1(66);
	sub_wire2(1, 67)    <= sub_wire1(67);
	sub_wire2(1, 68)    <= sub_wire1(68);
	sub_wire2(1, 69)    <= sub_wire1(69);
	sub_wire2(1, 70)    <= sub_wire1(70);
	sub_wire2(1, 71)    <= sub_wire1(71);
	sub_wire2(1, 72)    <= sub_wire1(72);
	sub_wire2(1, 73)    <= sub_wire1(73);
	sub_wire2(1, 74)    <= sub_wire1(74);
	sub_wire2(1, 75)    <= sub_wire1(75);
	sub_wire2(1, 76)    <= sub_wire1(76);
	sub_wire2(1, 77)    <= sub_wire1(77);
	sub_wire2(1, 78)    <= sub_wire1(78);
	sub_wire2(1, 79)    <= sub_wire1(79);
	sub_wire2(1, 80)    <= sub_wire1(80);
	sub_wire2(1, 81)    <= sub_wire1(81);
	sub_wire2(1, 82)    <= sub_wire1(82);
	sub_wire2(1, 83)    <= sub_wire1(83);
	sub_wire2(1, 84)    <= sub_wire1(84);
	sub_wire2(1, 85)    <= sub_wire1(85);
	sub_wire2(1, 86)    <= sub_wire1(86);
	sub_wire2(1, 87)    <= sub_wire1(87);
	sub_wire2(1, 88)    <= sub_wire1(88);
	sub_wire2(1, 89)    <= sub_wire1(89);
	sub_wire2(1, 90)    <= sub_wire1(90);
	sub_wire2(1, 91)    <= sub_wire1(91);
	sub_wire2(1, 92)    <= sub_wire1(92);
	sub_wire2(1, 93)    <= sub_wire1(93);
	sub_wire2(1, 94)    <= sub_wire1(94);
	sub_wire2(1, 95)    <= sub_wire1(95);
	sub_wire2(1, 96)    <= sub_wire1(96);
	sub_wire2(1, 97)    <= sub_wire1(97);
	sub_wire2(1, 98)    <= sub_wire1(98);
	sub_wire2(1, 99)    <= sub_wire1(99);
	sub_wire2(1, 100)    <= sub_wire1(100);
	sub_wire2(1, 101)    <= sub_wire1(101);
	sub_wire2(1, 102)    <= sub_wire1(102);
	sub_wire2(1, 103)    <= sub_wire1(103);
	sub_wire2(1, 104)    <= sub_wire1(104);
	sub_wire2(1, 105)    <= sub_wire1(105);
	sub_wire2(1, 106)    <= sub_wire1(106);
	sub_wire2(1, 107)    <= sub_wire1(107);
	sub_wire2(1, 108)    <= sub_wire1(108);
	sub_wire2(1, 109)    <= sub_wire1(109);
	sub_wire2(1, 110)    <= sub_wire1(110);
	sub_wire2(1, 111)    <= sub_wire1(111);
	sub_wire2(1, 112)    <= sub_wire1(112);
	sub_wire2(1, 113)    <= sub_wire1(113);
	sub_wire2(1, 114)    <= sub_wire1(114);
	sub_wire2(1, 115)    <= sub_wire1(115);
	sub_wire2(1, 116)    <= sub_wire1(116);
	sub_wire2(1, 117)    <= sub_wire1(117);
	sub_wire2(1, 118)    <= sub_wire1(118);
	sub_wire2(1, 119)    <= sub_wire1(119);
	sub_wire2(1, 120)    <= sub_wire1(120);
	sub_wire2(1, 121)    <= sub_wire1(121);
	sub_wire2(1, 122)    <= sub_wire1(122);
	sub_wire2(1, 123)    <= sub_wire1(123);
	sub_wire2(1, 124)    <= sub_wire1(124);
	sub_wire2(1, 125)    <= sub_wire1(125);
	sub_wire2(1, 126)    <= sub_wire1(126);
	sub_wire2(1, 127)    <= sub_wire1(127);
	sub_wire2(1, 128)    <= sub_wire1(128);
	sub_wire2(1, 129)    <= sub_wire1(129);
	sub_wire2(1, 130)    <= sub_wire1(130);
	sub_wire2(1, 131)    <= sub_wire1(131);
	sub_wire2(1, 132)    <= sub_wire1(132);
	sub_wire2(1, 133)    <= sub_wire1(133);
	sub_wire2(1, 134)    <= sub_wire1(134);
	sub_wire2(1, 135)    <= sub_wire1(135);
	sub_wire2(1, 136)    <= sub_wire1(136);
	sub_wire2(1, 137)    <= sub_wire1(137);
	sub_wire2(1, 138)    <= sub_wire1(138);
	sub_wire2(1, 139)    <= sub_wire1(139);
	sub_wire2(1, 140)    <= sub_wire1(140);
	sub_wire2(1, 141)    <= sub_wire1(141);
	sub_wire2(1, 142)    <= sub_wire1(142);
	sub_wire2(1, 143)    <= sub_wire1(143);
	sub_wire2(1, 144)    <= sub_wire1(144);
	sub_wire2(1, 145)    <= sub_wire1(145);
	sub_wire2(1, 146)    <= sub_wire1(146);
	sub_wire2(1, 147)    <= sub_wire1(147);
	sub_wire2(1, 148)    <= sub_wire1(148);
	sub_wire2(1, 149)    <= sub_wire1(149);
	sub_wire2(1, 150)    <= sub_wire1(150);
	sub_wire2(1, 151)    <= sub_wire1(151);
	sub_wire2(1, 152)    <= sub_wire1(152);
	sub_wire2(1, 153)    <= sub_wire1(153);
	sub_wire2(1, 154)    <= sub_wire1(154);
	sub_wire2(1, 155)    <= sub_wire1(155);
	sub_wire2(1, 156)    <= sub_wire1(156);
	sub_wire2(1, 157)    <= sub_wire1(157);
	sub_wire2(1, 158)    <= sub_wire1(158);
	sub_wire2(1, 159)    <= sub_wire1(159);
	sub_wire2(1, 160)    <= sub_wire1(160);
	sub_wire2(1, 161)    <= sub_wire1(161);
	sub_wire2(1, 162)    <= sub_wire1(162);
	sub_wire2(1, 163)    <= sub_wire1(163);
	sub_wire2(1, 164)    <= sub_wire1(164);
	sub_wire2(1, 165)    <= sub_wire1(165);
	sub_wire2(1, 166)    <= sub_wire1(166);
	sub_wire2(1, 167)    <= sub_wire1(167);
	sub_wire2(1, 168)    <= sub_wire1(168);
	sub_wire2(1, 169)    <= sub_wire1(169);
	sub_wire2(1, 170)    <= sub_wire1(170);
	sub_wire2(1, 171)    <= sub_wire1(171);
	sub_wire2(1, 172)    <= sub_wire1(172);
	sub_wire2(1, 173)    <= sub_wire1(173);
	sub_wire2(1, 174)    <= sub_wire1(174);
	sub_wire2(1, 175)    <= sub_wire1(175);
	sub_wire2(1, 176)    <= sub_wire1(176);
	sub_wire2(1, 177)    <= sub_wire1(177);
	sub_wire2(1, 178)    <= sub_wire1(178);
	sub_wire2(1, 179)    <= sub_wire1(179);
	sub_wire2(1, 180)    <= sub_wire1(180);
	sub_wire2(1, 181)    <= sub_wire1(181);
	sub_wire2(1, 182)    <= sub_wire1(182);
	sub_wire2(1, 183)    <= sub_wire1(183);
	sub_wire2(1, 184)    <= sub_wire1(184);
	sub_wire2(1, 185)    <= sub_wire1(185);
	sub_wire2(1, 186)    <= sub_wire1(186);
	sub_wire2(1, 187)    <= sub_wire1(187);
	sub_wire2(1, 188)    <= sub_wire1(188);
	sub_wire2(1, 189)    <= sub_wire1(189);
	sub_wire2(1, 190)    <= sub_wire1(190);
	sub_wire2(1, 191)    <= sub_wire1(191);
	sub_wire2(1, 192)    <= sub_wire1(192);
	sub_wire2(1, 193)    <= sub_wire1(193);
	sub_wire2(1, 194)    <= sub_wire1(194);
	sub_wire2(1, 195)    <= sub_wire1(195);
	sub_wire2(1, 196)    <= sub_wire1(196);
	sub_wire2(1, 197)    <= sub_wire1(197);
	sub_wire2(1, 198)    <= sub_wire1(198);
	sub_wire2(1, 199)    <= sub_wire1(199);
	sub_wire2(1, 200)    <= sub_wire1(200);
	sub_wire2(1, 201)    <= sub_wire1(201);
	sub_wire2(1, 202)    <= sub_wire1(202);
	sub_wire2(1, 203)    <= sub_wire1(203);
	sub_wire2(1, 204)    <= sub_wire1(204);
	sub_wire2(1, 205)    <= sub_wire1(205);
	sub_wire2(1, 206)    <= sub_wire1(206);
	sub_wire2(1, 207)    <= sub_wire1(207);
	sub_wire2(1, 208)    <= sub_wire1(208);
	sub_wire2(1, 209)    <= sub_wire1(209);
	sub_wire2(1, 210)    <= sub_wire1(210);
	sub_wire2(1, 211)    <= sub_wire1(211);
	sub_wire2(1, 212)    <= sub_wire1(212);
	sub_wire2(1, 213)    <= sub_wire1(213);
	sub_wire2(1, 214)    <= sub_wire1(214);
	sub_wire2(1, 215)    <= sub_wire1(215);
	sub_wire2(1, 216)    <= sub_wire1(216);
	sub_wire2(1, 217)    <= sub_wire1(217);
	sub_wire2(1, 218)    <= sub_wire1(218);
	sub_wire2(1, 219)    <= sub_wire1(219);
	sub_wire2(1, 220)    <= sub_wire1(220);
	sub_wire2(1, 221)    <= sub_wire1(221);
	sub_wire2(1, 222)    <= sub_wire1(222);
	sub_wire2(1, 223)    <= sub_wire1(223);
	sub_wire2(1, 224)    <= sub_wire1(224);
	sub_wire2(1, 225)    <= sub_wire1(225);
	sub_wire2(1, 226)    <= sub_wire1(226);
	sub_wire2(1, 227)    <= sub_wire1(227);
	sub_wire2(1, 228)    <= sub_wire1(228);
	sub_wire2(1, 229)    <= sub_wire1(229);
	sub_wire2(1, 230)    <= sub_wire1(230);
	sub_wire2(1, 231)    <= sub_wire1(231);
	sub_wire2(1, 232)    <= sub_wire1(232);
	sub_wire2(1, 233)    <= sub_wire1(233);
	sub_wire2(1, 234)    <= sub_wire1(234);
	sub_wire2(1, 235)    <= sub_wire1(235);
	sub_wire2(1, 236)    <= sub_wire1(236);
	sub_wire2(1, 237)    <= sub_wire1(237);
	sub_wire2(1, 238)    <= sub_wire1(238);
	sub_wire2(1, 239)    <= sub_wire1(239);
	sub_wire2(1, 240)    <= sub_wire1(240);
	sub_wire2(1, 241)    <= sub_wire1(241);
	sub_wire2(1, 242)    <= sub_wire1(242);
	sub_wire2(1, 243)    <= sub_wire1(243);
	sub_wire2(1, 244)    <= sub_wire1(244);
	sub_wire2(1, 245)    <= sub_wire1(245);
	sub_wire2(1, 246)    <= sub_wire1(246);
	sub_wire2(1, 247)    <= sub_wire1(247);
	sub_wire2(1, 248)    <= sub_wire1(248);
	sub_wire2(1, 249)    <= sub_wire1(249);
	sub_wire2(1, 250)    <= sub_wire1(250);
	sub_wire2(1, 251)    <= sub_wire1(251);
	sub_wire2(1, 252)    <= sub_wire1(252);
	sub_wire2(1, 253)    <= sub_wire1(253);
	sub_wire2(1, 254)    <= sub_wire1(254);
	sub_wire2(1, 255)    <= sub_wire1(255);
	sub_wire2(0, 0)    <= sub_wire3(0);
	sub_wire2(0, 1)    <= sub_wire3(1);
	sub_wire2(0, 2)    <= sub_wire3(2);
	sub_wire2(0, 3)    <= sub_wire3(3);
	sub_wire2(0, 4)    <= sub_wire3(4);
	sub_wire2(0, 5)    <= sub_wire3(5);
	sub_wire2(0, 6)    <= sub_wire3(6);
	sub_wire2(0, 7)    <= sub_wire3(7);
	sub_wire2(0, 8)    <= sub_wire3(8);
	sub_wire2(0, 9)    <= sub_wire3(9);
	sub_wire2(0, 10)    <= sub_wire3(10);
	sub_wire2(0, 11)    <= sub_wire3(11);
	sub_wire2(0, 12)    <= sub_wire3(12);
	sub_wire2(0, 13)    <= sub_wire3(13);
	sub_wire2(0, 14)    <= sub_wire3(14);
	sub_wire2(0, 15)    <= sub_wire3(15);
	sub_wire2(0, 16)    <= sub_wire3(16);
	sub_wire2(0, 17)    <= sub_wire3(17);
	sub_wire2(0, 18)    <= sub_wire3(18);
	sub_wire2(0, 19)    <= sub_wire3(19);
	sub_wire2(0, 20)    <= sub_wire3(20);
	sub_wire2(0, 21)    <= sub_wire3(21);
	sub_wire2(0, 22)    <= sub_wire3(22);
	sub_wire2(0, 23)    <= sub_wire3(23);
	sub_wire2(0, 24)    <= sub_wire3(24);
	sub_wire2(0, 25)    <= sub_wire3(25);
	sub_wire2(0, 26)    <= sub_wire3(26);
	sub_wire2(0, 27)    <= sub_wire3(27);
	sub_wire2(0, 28)    <= sub_wire3(28);
	sub_wire2(0, 29)    <= sub_wire3(29);
	sub_wire2(0, 30)    <= sub_wire3(30);
	sub_wire2(0, 31)    <= sub_wire3(31);
	sub_wire2(0, 32)    <= sub_wire3(32);
	sub_wire2(0, 33)    <= sub_wire3(33);
	sub_wire2(0, 34)    <= sub_wire3(34);
	sub_wire2(0, 35)    <= sub_wire3(35);
	sub_wire2(0, 36)    <= sub_wire3(36);
	sub_wire2(0, 37)    <= sub_wire3(37);
	sub_wire2(0, 38)    <= sub_wire3(38);
	sub_wire2(0, 39)    <= sub_wire3(39);
	sub_wire2(0, 40)    <= sub_wire3(40);
	sub_wire2(0, 41)    <= sub_wire3(41);
	sub_wire2(0, 42)    <= sub_wire3(42);
	sub_wire2(0, 43)    <= sub_wire3(43);
	sub_wire2(0, 44)    <= sub_wire3(44);
	sub_wire2(0, 45)    <= sub_wire3(45);
	sub_wire2(0, 46)    <= sub_wire3(46);
	sub_wire2(0, 47)    <= sub_wire3(47);
	sub_wire2(0, 48)    <= sub_wire3(48);
	sub_wire2(0, 49)    <= sub_wire3(49);
	sub_wire2(0, 50)    <= sub_wire3(50);
	sub_wire2(0, 51)    <= sub_wire3(51);
	sub_wire2(0, 52)    <= sub_wire3(52);
	sub_wire2(0, 53)    <= sub_wire3(53);
	sub_wire2(0, 54)    <= sub_wire3(54);
	sub_wire2(0, 55)    <= sub_wire3(55);
	sub_wire2(0, 56)    <= sub_wire3(56);
	sub_wire2(0, 57)    <= sub_wire3(57);
	sub_wire2(0, 58)    <= sub_wire3(58);
	sub_wire2(0, 59)    <= sub_wire3(59);
	sub_wire2(0, 60)    <= sub_wire3(60);
	sub_wire2(0, 61)    <= sub_wire3(61);
	sub_wire2(0, 62)    <= sub_wire3(62);
	sub_wire2(0, 63)    <= sub_wire3(63);
	sub_wire2(0, 64)    <= sub_wire3(64);
	sub_wire2(0, 65)    <= sub_wire3(65);
	sub_wire2(0, 66)    <= sub_wire3(66);
	sub_wire2(0, 67)    <= sub_wire3(67);
	sub_wire2(0, 68)    <= sub_wire3(68);
	sub_wire2(0, 69)    <= sub_wire3(69);
	sub_wire2(0, 70)    <= sub_wire3(70);
	sub_wire2(0, 71)    <= sub_wire3(71);
	sub_wire2(0, 72)    <= sub_wire3(72);
	sub_wire2(0, 73)    <= sub_wire3(73);
	sub_wire2(0, 74)    <= sub_wire3(74);
	sub_wire2(0, 75)    <= sub_wire3(75);
	sub_wire2(0, 76)    <= sub_wire3(76);
	sub_wire2(0, 77)    <= sub_wire3(77);
	sub_wire2(0, 78)    <= sub_wire3(78);
	sub_wire2(0, 79)    <= sub_wire3(79);
	sub_wire2(0, 80)    <= sub_wire3(80);
	sub_wire2(0, 81)    <= sub_wire3(81);
	sub_wire2(0, 82)    <= sub_wire3(82);
	sub_wire2(0, 83)    <= sub_wire3(83);
	sub_wire2(0, 84)    <= sub_wire3(84);
	sub_wire2(0, 85)    <= sub_wire3(85);
	sub_wire2(0, 86)    <= sub_wire3(86);
	sub_wire2(0, 87)    <= sub_wire3(87);
	sub_wire2(0, 88)    <= sub_wire3(88);
	sub_wire2(0, 89)    <= sub_wire3(89);
	sub_wire2(0, 90)    <= sub_wire3(90);
	sub_wire2(0, 91)    <= sub_wire3(91);
	sub_wire2(0, 92)    <= sub_wire3(92);
	sub_wire2(0, 93)    <= sub_wire3(93);
	sub_wire2(0, 94)    <= sub_wire3(94);
	sub_wire2(0, 95)    <= sub_wire3(95);
	sub_wire2(0, 96)    <= sub_wire3(96);
	sub_wire2(0, 97)    <= sub_wire3(97);
	sub_wire2(0, 98)    <= sub_wire3(98);
	sub_wire2(0, 99)    <= sub_wire3(99);
	sub_wire2(0, 100)    <= sub_wire3(100);
	sub_wire2(0, 101)    <= sub_wire3(101);
	sub_wire2(0, 102)    <= sub_wire3(102);
	sub_wire2(0, 103)    <= sub_wire3(103);
	sub_wire2(0, 104)    <= sub_wire3(104);
	sub_wire2(0, 105)    <= sub_wire3(105);
	sub_wire2(0, 106)    <= sub_wire3(106);
	sub_wire2(0, 107)    <= sub_wire3(107);
	sub_wire2(0, 108)    <= sub_wire3(108);
	sub_wire2(0, 109)    <= sub_wire3(109);
	sub_wire2(0, 110)    <= sub_wire3(110);
	sub_wire2(0, 111)    <= sub_wire3(111);
	sub_wire2(0, 112)    <= sub_wire3(112);
	sub_wire2(0, 113)    <= sub_wire3(113);
	sub_wire2(0, 114)    <= sub_wire3(114);
	sub_wire2(0, 115)    <= sub_wire3(115);
	sub_wire2(0, 116)    <= sub_wire3(116);
	sub_wire2(0, 117)    <= sub_wire3(117);
	sub_wire2(0, 118)    <= sub_wire3(118);
	sub_wire2(0, 119)    <= sub_wire3(119);
	sub_wire2(0, 120)    <= sub_wire3(120);
	sub_wire2(0, 121)    <= sub_wire3(121);
	sub_wire2(0, 122)    <= sub_wire3(122);
	sub_wire2(0, 123)    <= sub_wire3(123);
	sub_wire2(0, 124)    <= sub_wire3(124);
	sub_wire2(0, 125)    <= sub_wire3(125);
	sub_wire2(0, 126)    <= sub_wire3(126);
	sub_wire2(0, 127)    <= sub_wire3(127);
	sub_wire2(0, 128)    <= sub_wire3(128);
	sub_wire2(0, 129)    <= sub_wire3(129);
	sub_wire2(0, 130)    <= sub_wire3(130);
	sub_wire2(0, 131)    <= sub_wire3(131);
	sub_wire2(0, 132)    <= sub_wire3(132);
	sub_wire2(0, 133)    <= sub_wire3(133);
	sub_wire2(0, 134)    <= sub_wire3(134);
	sub_wire2(0, 135)    <= sub_wire3(135);
	sub_wire2(0, 136)    <= sub_wire3(136);
	sub_wire2(0, 137)    <= sub_wire3(137);
	sub_wire2(0, 138)    <= sub_wire3(138);
	sub_wire2(0, 139)    <= sub_wire3(139);
	sub_wire2(0, 140)    <= sub_wire3(140);
	sub_wire2(0, 141)    <= sub_wire3(141);
	sub_wire2(0, 142)    <= sub_wire3(142);
	sub_wire2(0, 143)    <= sub_wire3(143);
	sub_wire2(0, 144)    <= sub_wire3(144);
	sub_wire2(0, 145)    <= sub_wire3(145);
	sub_wire2(0, 146)    <= sub_wire3(146);
	sub_wire2(0, 147)    <= sub_wire3(147);
	sub_wire2(0, 148)    <= sub_wire3(148);
	sub_wire2(0, 149)    <= sub_wire3(149);
	sub_wire2(0, 150)    <= sub_wire3(150);
	sub_wire2(0, 151)    <= sub_wire3(151);
	sub_wire2(0, 152)    <= sub_wire3(152);
	sub_wire2(0, 153)    <= sub_wire3(153);
	sub_wire2(0, 154)    <= sub_wire3(154);
	sub_wire2(0, 155)    <= sub_wire3(155);
	sub_wire2(0, 156)    <= sub_wire3(156);
	sub_wire2(0, 157)    <= sub_wire3(157);
	sub_wire2(0, 158)    <= sub_wire3(158);
	sub_wire2(0, 159)    <= sub_wire3(159);
	sub_wire2(0, 160)    <= sub_wire3(160);
	sub_wire2(0, 161)    <= sub_wire3(161);
	sub_wire2(0, 162)    <= sub_wire3(162);
	sub_wire2(0, 163)    <= sub_wire3(163);
	sub_wire2(0, 164)    <= sub_wire3(164);
	sub_wire2(0, 165)    <= sub_wire3(165);
	sub_wire2(0, 166)    <= sub_wire3(166);
	sub_wire2(0, 167)    <= sub_wire3(167);
	sub_wire2(0, 168)    <= sub_wire3(168);
	sub_wire2(0, 169)    <= sub_wire3(169);
	sub_wire2(0, 170)    <= sub_wire3(170);
	sub_wire2(0, 171)    <= sub_wire3(171);
	sub_wire2(0, 172)    <= sub_wire3(172);
	sub_wire2(0, 173)    <= sub_wire3(173);
	sub_wire2(0, 174)    <= sub_wire3(174);
	sub_wire2(0, 175)    <= sub_wire3(175);
	sub_wire2(0, 176)    <= sub_wire3(176);
	sub_wire2(0, 177)    <= sub_wire3(177);
	sub_wire2(0, 178)    <= sub_wire3(178);
	sub_wire2(0, 179)    <= sub_wire3(179);
	sub_wire2(0, 180)    <= sub_wire3(180);
	sub_wire2(0, 181)    <= sub_wire3(181);
	sub_wire2(0, 182)    <= sub_wire3(182);
	sub_wire2(0, 183)    <= sub_wire3(183);
	sub_wire2(0, 184)    <= sub_wire3(184);
	sub_wire2(0, 185)    <= sub_wire3(185);
	sub_wire2(0, 186)    <= sub_wire3(186);
	sub_wire2(0, 187)    <= sub_wire3(187);
	sub_wire2(0, 188)    <= sub_wire3(188);
	sub_wire2(0, 189)    <= sub_wire3(189);
	sub_wire2(0, 190)    <= sub_wire3(190);
	sub_wire2(0, 191)    <= sub_wire3(191);
	sub_wire2(0, 192)    <= sub_wire3(192);
	sub_wire2(0, 193)    <= sub_wire3(193);
	sub_wire2(0, 194)    <= sub_wire3(194);
	sub_wire2(0, 195)    <= sub_wire3(195);
	sub_wire2(0, 196)    <= sub_wire3(196);
	sub_wire2(0, 197)    <= sub_wire3(197);
	sub_wire2(0, 198)    <= sub_wire3(198);
	sub_wire2(0, 199)    <= sub_wire3(199);
	sub_wire2(0, 200)    <= sub_wire3(200);
	sub_wire2(0, 201)    <= sub_wire3(201);
	sub_wire2(0, 202)    <= sub_wire3(202);
	sub_wire2(0, 203)    <= sub_wire3(203);
	sub_wire2(0, 204)    <= sub_wire3(204);
	sub_wire2(0, 205)    <= sub_wire3(205);
	sub_wire2(0, 206)    <= sub_wire3(206);
	sub_wire2(0, 207)    <= sub_wire3(207);
	sub_wire2(0, 208)    <= sub_wire3(208);
	sub_wire2(0, 209)    <= sub_wire3(209);
	sub_wire2(0, 210)    <= sub_wire3(210);
	sub_wire2(0, 211)    <= sub_wire3(211);
	sub_wire2(0, 212)    <= sub_wire3(212);
	sub_wire2(0, 213)    <= sub_wire3(213);
	sub_wire2(0, 214)    <= sub_wire3(214);
	sub_wire2(0, 215)    <= sub_wire3(215);
	sub_wire2(0, 216)    <= sub_wire3(216);
	sub_wire2(0, 217)    <= sub_wire3(217);
	sub_wire2(0, 218)    <= sub_wire3(218);
	sub_wire2(0, 219)    <= sub_wire3(219);
	sub_wire2(0, 220)    <= sub_wire3(220);
	sub_wire2(0, 221)    <= sub_wire3(221);
	sub_wire2(0, 222)    <= sub_wire3(222);
	sub_wire2(0, 223)    <= sub_wire3(223);
	sub_wire2(0, 224)    <= sub_wire3(224);
	sub_wire2(0, 225)    <= sub_wire3(225);
	sub_wire2(0, 226)    <= sub_wire3(226);
	sub_wire2(0, 227)    <= sub_wire3(227);
	sub_wire2(0, 228)    <= sub_wire3(228);
	sub_wire2(0, 229)    <= sub_wire3(229);
	sub_wire2(0, 230)    <= sub_wire3(230);
	sub_wire2(0, 231)    <= sub_wire3(231);
	sub_wire2(0, 232)    <= sub_wire3(232);
	sub_wire2(0, 233)    <= sub_wire3(233);
	sub_wire2(0, 234)    <= sub_wire3(234);
	sub_wire2(0, 235)    <= sub_wire3(235);
	sub_wire2(0, 236)    <= sub_wire3(236);
	sub_wire2(0, 237)    <= sub_wire3(237);
	sub_wire2(0, 238)    <= sub_wire3(238);
	sub_wire2(0, 239)    <= sub_wire3(239);
	sub_wire2(0, 240)    <= sub_wire3(240);
	sub_wire2(0, 241)    <= sub_wire3(241);
	sub_wire2(0, 242)    <= sub_wire3(242);
	sub_wire2(0, 243)    <= sub_wire3(243);
	sub_wire2(0, 244)    <= sub_wire3(244);
	sub_wire2(0, 245)    <= sub_wire3(245);
	sub_wire2(0, 246)    <= sub_wire3(246);
	sub_wire2(0, 247)    <= sub_wire3(247);
	sub_wire2(0, 248)    <= sub_wire3(248);
	sub_wire2(0, 249)    <= sub_wire3(249);
	sub_wire2(0, 250)    <= sub_wire3(250);
	sub_wire2(0, 251)    <= sub_wire3(251);
	sub_wire2(0, 252)    <= sub_wire3(252);
	sub_wire2(0, 253)    <= sub_wire3(253);
	sub_wire2(0, 254)    <= sub_wire3(254);
	sub_wire2(0, 255)    <= sub_wire3(255);
	sub_wire4    <= sel;
	sub_wire5(0)    <= sub_wire4;

	LPM_MUX_component : LPM_MUX
	GENERIC MAP (
		lpm_size => 2,
		lpm_type => "LPM_MUX",
		lpm_width => 256,
		lpm_widths => 1
	)
	PORT MAP (
		data => sub_wire2,
		sel => sub_wire5,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "2"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "256"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "1"
-- Retrieval info: USED_PORT: data0x 0 0 256 0 INPUT NODEFVAL "data0x[255..0]"
-- Retrieval info: USED_PORT: data1x 0 0 256 0 INPUT NODEFVAL "data1x[255..0]"
-- Retrieval info: USED_PORT: result 0 0 256 0 OUTPUT NODEFVAL "result[255..0]"
-- Retrieval info: USED_PORT: sel 0 0 0 0 INPUT NODEFVAL "sel"
-- Retrieval info: CONNECT: @data 1 0 256 0 data0x 0 0 256 0
-- Retrieval info: CONNECT: @data 1 1 256 0 data1x 0 0 256 0
-- Retrieval info: CONNECT: @sel 0 0 1 0 sel 0 0 0 0
-- Retrieval info: CONNECT: result 0 0 256 0 @result 0 0 256 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux256.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux256.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux256.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux256.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux256_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
