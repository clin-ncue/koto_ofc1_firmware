// megafunction wizard: %PARALLEL_ADD%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: parallel_add 

// ============================================================
// File Name: parallel_add37_8b.v
// Megafunction Name(s):
// 			parallel_add
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 15.0.0 Build 145 04/22/2015 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, the Altera Quartus II License Agreement,
//the Altera MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Altera and sold by Altera or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module parallel_add37_8b (
	clock,
	data0x,
	data10x,
	data11x,
	data12x,
	data13x,
	data14x,
	data15x,
	data16x,
	data17x,
	data18x,
	data19x,
	data1x,
	data20x,
	data21x,
	data22x,
	data23x,
	data24x,
	data25x,
	data26x,
	data27x,
	data28x,
	data29x,
	data2x,
	data30x,
	data31x,
	data32x,
	data33x,
	data34x,
	data35x,
	data36x,
	data3x,
	data4x,
	data5x,
	data6x,
	data7x,
	data8x,
	data9x,
	result);

	input	  clock;
	input	[7:0]  data0x;
	input	[7:0]  data10x;
	input	[7:0]  data11x;
	input	[7:0]  data12x;
	input	[7:0]  data13x;
	input	[7:0]  data14x;
	input	[7:0]  data15x;
	input	[7:0]  data16x;
	input	[7:0]  data17x;
	input	[7:0]  data18x;
	input	[7:0]  data19x;
	input	[7:0]  data1x;
	input	[7:0]  data20x;
	input	[7:0]  data21x;
	input	[7:0]  data22x;
	input	[7:0]  data23x;
	input	[7:0]  data24x;
	input	[7:0]  data25x;
	input	[7:0]  data26x;
	input	[7:0]  data27x;
	input	[7:0]  data28x;
	input	[7:0]  data29x;
	input	[7:0]  data2x;
	input	[7:0]  data30x;
	input	[7:0]  data31x;
	input	[7:0]  data32x;
	input	[7:0]  data33x;
	input	[7:0]  data34x;
	input	[7:0]  data35x;
	input	[7:0]  data36x;
	input	[7:0]  data3x;
	input	[7:0]  data4x;
	input	[7:0]  data5x;
	input	[7:0]  data6x;
	input	[7:0]  data7x;
	input	[7:0]  data8x;
	input	[7:0]  data9x;
	output	[13:0]  result;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri0	  clock;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [13:0] sub_wire38;
	wire [7:0] sub_wire37 = data36x[7:0];
	wire [7:0] sub_wire36 = data35x[7:0];
	wire [7:0] sub_wire35 = data34x[7:0];
	wire [7:0] sub_wire34 = data33x[7:0];
	wire [7:0] sub_wire33 = data32x[7:0];
	wire [7:0] sub_wire32 = data31x[7:0];
	wire [7:0] sub_wire31 = data30x[7:0];
	wire [7:0] sub_wire30 = data29x[7:0];
	wire [7:0] sub_wire29 = data28x[7:0];
	wire [7:0] sub_wire28 = data27x[7:0];
	wire [7:0] sub_wire27 = data26x[7:0];
	wire [7:0] sub_wire26 = data25x[7:0];
	wire [7:0] sub_wire25 = data24x[7:0];
	wire [7:0] sub_wire24 = data23x[7:0];
	wire [7:0] sub_wire23 = data22x[7:0];
	wire [7:0] sub_wire22 = data21x[7:0];
	wire [7:0] sub_wire21 = data20x[7:0];
	wire [7:0] sub_wire20 = data19x[7:0];
	wire [7:0] sub_wire19 = data18x[7:0];
	wire [7:0] sub_wire18 = data17x[7:0];
	wire [7:0] sub_wire17 = data16x[7:0];
	wire [7:0] sub_wire16 = data15x[7:0];
	wire [7:0] sub_wire15 = data14x[7:0];
	wire [7:0] sub_wire14 = data13x[7:0];
	wire [7:0] sub_wire13 = data12x[7:0];
	wire [7:0] sub_wire12 = data11x[7:0];
	wire [7:0] sub_wire11 = data10x[7:0];
	wire [7:0] sub_wire10 = data9x[7:0];
	wire [7:0] sub_wire9 = data8x[7:0];
	wire [7:0] sub_wire8 = data7x[7:0];
	wire [7:0] sub_wire7 = data6x[7:0];
	wire [7:0] sub_wire6 = data5x[7:0];
	wire [7:0] sub_wire5 = data4x[7:0];
	wire [7:0] sub_wire4 = data3x[7:0];
	wire [7:0] sub_wire3 = data2x[7:0];
	wire [7:0] sub_wire2 = data1x[7:0];
	wire [7:0] sub_wire0 = data0x[7:0];
	wire [295:0] sub_wire1 = {sub_wire37, sub_wire36, sub_wire35, sub_wire34, sub_wire33, sub_wire32, sub_wire31, sub_wire30, sub_wire29, sub_wire28, sub_wire27, sub_wire26, sub_wire25, sub_wire24, sub_wire23, sub_wire22, sub_wire21, sub_wire20, sub_wire19, sub_wire18, sub_wire17, sub_wire16, sub_wire15, sub_wire14, sub_wire13, sub_wire12, sub_wire11, sub_wire10, sub_wire9, sub_wire8, sub_wire7, sub_wire6, sub_wire5, sub_wire4, sub_wire3, sub_wire2, sub_wire0};
	wire [13:0] result = sub_wire38[13:0];

	parallel_add	parallel_add_component (
				.clock (clock),
				.data (sub_wire1),
				.result (sub_wire38)
				// synopsys translate_off
				,
				.aclr (),
				.clken ()
				// synopsys translate_on
				);
	defparam
		parallel_add_component.msw_subtract = "NO",
		parallel_add_component.pipeline = 1,
		parallel_add_component.representation = "UNSIGNED",
		parallel_add_component.result_alignment = "LSB",
		parallel_add_component.shift = 0,
		parallel_add_component.size = 37,
		parallel_add_component.width = 8,
		parallel_add_component.widthr = 14;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: MSW_SUBTRACT STRING "NO"
// Retrieval info: CONSTANT: PIPELINE NUMERIC "1"
// Retrieval info: CONSTANT: REPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: RESULT_ALIGNMENT STRING "LSB"
// Retrieval info: CONSTANT: SHIFT NUMERIC "0"
// Retrieval info: CONSTANT: SIZE NUMERIC "37"
// Retrieval info: CONSTANT: WIDTH NUMERIC "8"
// Retrieval info: CONSTANT: WIDTHR NUMERIC "14"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT GND "clock"
// Retrieval info: USED_PORT: data0x 0 0 8 0 INPUT NODEFVAL "data0x[7..0]"
// Retrieval info: USED_PORT: data10x 0 0 8 0 INPUT NODEFVAL "data10x[7..0]"
// Retrieval info: USED_PORT: data11x 0 0 8 0 INPUT NODEFVAL "data11x[7..0]"
// Retrieval info: USED_PORT: data12x 0 0 8 0 INPUT NODEFVAL "data12x[7..0]"
// Retrieval info: USED_PORT: data13x 0 0 8 0 INPUT NODEFVAL "data13x[7..0]"
// Retrieval info: USED_PORT: data14x 0 0 8 0 INPUT NODEFVAL "data14x[7..0]"
// Retrieval info: USED_PORT: data15x 0 0 8 0 INPUT NODEFVAL "data15x[7..0]"
// Retrieval info: USED_PORT: data16x 0 0 8 0 INPUT NODEFVAL "data16x[7..0]"
// Retrieval info: USED_PORT: data17x 0 0 8 0 INPUT NODEFVAL "data17x[7..0]"
// Retrieval info: USED_PORT: data18x 0 0 8 0 INPUT NODEFVAL "data18x[7..0]"
// Retrieval info: USED_PORT: data19x 0 0 8 0 INPUT NODEFVAL "data19x[7..0]"
// Retrieval info: USED_PORT: data1x 0 0 8 0 INPUT NODEFVAL "data1x[7..0]"
// Retrieval info: USED_PORT: data20x 0 0 8 0 INPUT NODEFVAL "data20x[7..0]"
// Retrieval info: USED_PORT: data21x 0 0 8 0 INPUT NODEFVAL "data21x[7..0]"
// Retrieval info: USED_PORT: data22x 0 0 8 0 INPUT NODEFVAL "data22x[7..0]"
// Retrieval info: USED_PORT: data23x 0 0 8 0 INPUT NODEFVAL "data23x[7..0]"
// Retrieval info: USED_PORT: data24x 0 0 8 0 INPUT NODEFVAL "data24x[7..0]"
// Retrieval info: USED_PORT: data25x 0 0 8 0 INPUT NODEFVAL "data25x[7..0]"
// Retrieval info: USED_PORT: data26x 0 0 8 0 INPUT NODEFVAL "data26x[7..0]"
// Retrieval info: USED_PORT: data27x 0 0 8 0 INPUT NODEFVAL "data27x[7..0]"
// Retrieval info: USED_PORT: data28x 0 0 8 0 INPUT NODEFVAL "data28x[7..0]"
// Retrieval info: USED_PORT: data29x 0 0 8 0 INPUT NODEFVAL "data29x[7..0]"
// Retrieval info: USED_PORT: data2x 0 0 8 0 INPUT NODEFVAL "data2x[7..0]"
// Retrieval info: USED_PORT: data30x 0 0 8 0 INPUT NODEFVAL "data30x[7..0]"
// Retrieval info: USED_PORT: data31x 0 0 8 0 INPUT NODEFVAL "data31x[7..0]"
// Retrieval info: USED_PORT: data32x 0 0 8 0 INPUT NODEFVAL "data32x[7..0]"
// Retrieval info: USED_PORT: data33x 0 0 8 0 INPUT NODEFVAL "data33x[7..0]"
// Retrieval info: USED_PORT: data34x 0 0 8 0 INPUT NODEFVAL "data34x[7..0]"
// Retrieval info: USED_PORT: data35x 0 0 8 0 INPUT NODEFVAL "data35x[7..0]"
// Retrieval info: USED_PORT: data36x 0 0 8 0 INPUT NODEFVAL "data36x[7..0]"
// Retrieval info: USED_PORT: data3x 0 0 8 0 INPUT NODEFVAL "data3x[7..0]"
// Retrieval info: USED_PORT: data4x 0 0 8 0 INPUT NODEFVAL "data4x[7..0]"
// Retrieval info: USED_PORT: data5x 0 0 8 0 INPUT NODEFVAL "data5x[7..0]"
// Retrieval info: USED_PORT: data6x 0 0 8 0 INPUT NODEFVAL "data6x[7..0]"
// Retrieval info: USED_PORT: data7x 0 0 8 0 INPUT NODEFVAL "data7x[7..0]"
// Retrieval info: USED_PORT: data8x 0 0 8 0 INPUT NODEFVAL "data8x[7..0]"
// Retrieval info: USED_PORT: data9x 0 0 8 0 INPUT NODEFVAL "data9x[7..0]"
// Retrieval info: USED_PORT: result 0 0 14 0 OUTPUT NODEFVAL "result[13..0]"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 8 0 data0x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 80 data10x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 88 data11x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 96 data12x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 104 data13x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 112 data14x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 120 data15x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 128 data16x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 136 data17x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 144 data18x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 152 data19x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 8 data1x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 160 data20x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 168 data21x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 176 data22x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 184 data23x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 192 data24x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 200 data25x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 208 data26x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 216 data27x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 224 data28x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 232 data29x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 16 data2x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 240 data30x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 248 data31x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 256 data32x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 264 data33x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 272 data34x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 280 data35x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 288 data36x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 24 data3x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 32 data4x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 40 data5x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 48 data6x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 56 data7x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 64 data8x 0 0 8 0
// Retrieval info: CONNECT: @data 0 0 8 72 data9x 0 0 8 0
// Retrieval info: CONNECT: result 0 0 14 0 @result 0 0 14 0
// Retrieval info: GEN_FILE: TYPE_NORMAL parallel_add37_8b.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL parallel_add37_8b.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL parallel_add37_8b.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL parallel_add37_8b.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL parallel_add37_8b_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL parallel_add37_8b_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
